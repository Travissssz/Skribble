`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/11/2025 12:44:19 AM
// Design Name: 
// Module Name: timer_frame
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module timer_frame(input frame_rate, input [12:0] pixel_index, output reg [15:0] oled_data);
    reg [15:0] frame_count = 1;
    parameter picture_total_count = 1;
    
    always @ (posedge frame_rate) begin
        frame_count <= (frame_count == picture_total_count - 1) ? 0 : frame_count + 1;
    end
   
    always @ (*) begin
        if (((pixel_index >= 411) && (pixel_index <= 418)) || ((pixel_index >= 421) && (pixel_index <= 426)) || ((pixel_index >= 429) && (pixel_index <= 430)) || ((pixel_index >= 434) && (pixel_index <= 435)) || ((pixel_index >= 438) && (pixel_index <= 443)) || ((pixel_index >= 446) && (pixel_index <= 449)) || ((pixel_index >= 507) && (pixel_index <= 514)) || ((pixel_index >= 517) && (pixel_index <= 522)) || ((pixel_index >= 525) && (pixel_index <= 526)) || ((pixel_index >= 530) && (pixel_index <= 531)) || ((pixel_index >= 534) && (pixel_index <= 539)) || ((pixel_index >= 542) && (pixel_index <= 546)) || ((pixel_index >= 606) && (pixel_index <= 607)) || ((pixel_index >= 615) && (pixel_index <= 616)) || ((pixel_index >= 621) && (pixel_index <= 623)) || ((pixel_index >= 625) && (pixel_index <= 627)) || ((pixel_index >= 630) && (pixel_index <= 631)) || ((pixel_index >= 638) && (pixel_index <= 639)) || ((pixel_index >= 642) && (pixel_index <= 643)) || ((pixel_index >= 702) && (pixel_index <= 703)) || ((pixel_index >= 711) && (pixel_index <= 712)) || ((pixel_index >= 717) && (pixel_index <= 723)) || ((pixel_index >= 726) && (pixel_index <= 727)) || ((pixel_index >= 734) && (pixel_index <= 735)) || ((pixel_index >= 738) && (pixel_index <= 739)) || ((pixel_index >= 798) && (pixel_index <= 799)) || ((pixel_index >= 807) && (pixel_index <= 808)) || ((pixel_index >= 813) && (pixel_index <= 814)) || pixel_index == 816 || ((pixel_index >= 818) && (pixel_index <= 819)) || ((pixel_index >= 822) && (pixel_index <= 826)) || ((pixel_index >= 830) && (pixel_index <= 834)) || ((pixel_index >= 894) && (pixel_index <= 895)) || ((pixel_index >= 903) && (pixel_index <= 904)) || ((pixel_index >= 909) && (pixel_index <= 910)) || ((pixel_index >= 914) && (pixel_index <= 915)) || ((pixel_index >= 918) && (pixel_index <= 922)) || ((pixel_index >= 926) && (pixel_index <= 929)) || ((pixel_index >= 990) && (pixel_index <= 991)) || ((pixel_index >= 999) && (pixel_index <= 1000)) || ((pixel_index >= 1005) && (pixel_index <= 1006)) || ((pixel_index >= 1010) && (pixel_index <= 1011)) || ((pixel_index >= 1014) && (pixel_index <= 1015)) || ((pixel_index >= 1022) && (pixel_index <= 1024)) || ((pixel_index >= 1086) && (pixel_index <= 1087)) || ((pixel_index >= 1095) && (pixel_index <= 1096)) || ((pixel_index >= 1101) && (pixel_index <= 1102)) || ((pixel_index >= 1106) && (pixel_index <= 1107)) || ((pixel_index >= 1110) && (pixel_index <= 1111)) || ((pixel_index >= 1118) && (pixel_index <= 1122)) || ((pixel_index >= 1182) && (pixel_index <= 1183)) || ((pixel_index >= 1189) && (pixel_index <= 1194)) || ((pixel_index >= 1197) && (pixel_index <= 1198)) || ((pixel_index >= 1202) && (pixel_index <= 1203)) || ((pixel_index >= 1206) && (pixel_index <= 1211)) || ((pixel_index >= 1214) && (pixel_index <= 1215)) || ((pixel_index >= 1217) && (pixel_index <= 1219)) || ((pixel_index >= 1278) && (pixel_index <= 1279)) || ((pixel_index >= 1285) && (pixel_index <= 1290)) || ((pixel_index >= 1293) && (pixel_index <= 1294)) || ((pixel_index >= 1298) && (pixel_index <= 1299)) || ((pixel_index >= 1302) && (pixel_index <= 1307)) || ((pixel_index >= 1310) && (pixel_index <= 1311)) || ((pixel_index >= 1314) && (pixel_index <= 1315)) || ((pixel_index >= 2116) && (pixel_index <= 2134)) || ((pixel_index >= 2139) && (pixel_index <= 2157)) || ((pixel_index >= 2162) && (pixel_index <= 2180)) || ((pixel_index >= 2185) && (pixel_index <= 2203)) || pixel_index == 2212 || pixel_index == 2230 || pixel_index == 2235 || pixel_index == 2253 || pixel_index == 2258 || pixel_index == 2276 || pixel_index == 2281 || pixel_index == 2299 || pixel_index == 2308 || pixel_index == 2326 || pixel_index == 2331 || pixel_index == 2349 || pixel_index == 2354 || pixel_index == 2372 || pixel_index == 2377 || pixel_index == 2395 || pixel_index == 2404 || ((pixel_index >= 2410) && (pixel_index <= 2416)) || pixel_index == 2422 || pixel_index == 2427 || ((pixel_index >= 2433) && (pixel_index <= 2439)) || pixel_index == 2445 || pixel_index == 2450 || ((pixel_index >= 2458) && (pixel_index <= 2459)) || pixel_index == 2468 || pixel_index == 2473 || ((pixel_index >= 2479) && (pixel_index <= 2485)) || pixel_index == 2491 || pixel_index == 2500 || ((pixel_index >= 2506) && (pixel_index <= 2512)) || pixel_index == 2518 || pixel_index == 2523 || ((pixel_index >= 2529) && (pixel_index <= 2535)) || pixel_index == 2541 || pixel_index == 2546 || ((pixel_index >= 2554) && (pixel_index <= 2555)) || pixel_index == 2564 || pixel_index == 2569 || ((pixel_index >= 2575) && (pixel_index <= 2581)) || pixel_index == 2587 || pixel_index == 2596 || ((pixel_index >= 2607) && (pixel_index <= 2608)) || pixel_index == 2614 || pixel_index == 2619 || ((pixel_index >= 2630) && (pixel_index <= 2631)) || pixel_index == 2637 || pixel_index == 2642 || ((pixel_index >= 2650) && (pixel_index <= 2651)) || pixel_index == 2660 || pixel_index == 2665 || ((pixel_index >= 2671) && (pixel_index <= 2672)) || ((pixel_index >= 2676) && (pixel_index <= 2677)) || pixel_index == 2683 || pixel_index == 2692 || ((pixel_index >= 2703) && (pixel_index <= 2704)) || pixel_index == 2710 || pixel_index == 2715 || ((pixel_index >= 2726) && (pixel_index <= 2727)) || pixel_index == 2733 || pixel_index == 2738 || ((pixel_index >= 2746) && (pixel_index <= 2747)) || pixel_index == 2756 || pixel_index == 2761 || ((pixel_index >= 2767) && (pixel_index <= 2768)) || ((pixel_index >= 2772) && (pixel_index <= 2773)) || pixel_index == 2779 || pixel_index == 2788 || ((pixel_index >= 2799) && (pixel_index <= 2800)) || pixel_index == 2806 || pixel_index == 2811 || ((pixel_index >= 2822) && (pixel_index <= 2823)) || pixel_index == 2829 || pixel_index == 2834 || ((pixel_index >= 2842) && (pixel_index <= 2843)) || pixel_index == 2852 || pixel_index == 2857 || ((pixel_index >= 2863) && (pixel_index <= 2864)) || ((pixel_index >= 2868) && (pixel_index <= 2869)) || pixel_index == 2875 || pixel_index == 2884 || ((pixel_index >= 2890) && (pixel_index <= 2896)) || pixel_index == 2902 || pixel_index == 2907 || ((pixel_index >= 2913) && (pixel_index <= 2919)) || pixel_index == 2925 || pixel_index == 2930 || ((pixel_index >= 2938) && (pixel_index <= 2939)) || pixel_index == 2948 || pixel_index == 2953 || ((pixel_index >= 2959) && (pixel_index <= 2960)) || ((pixel_index >= 2964) && (pixel_index <= 2965)) || pixel_index == 2971 || pixel_index == 2980 || ((pixel_index >= 2986) && (pixel_index <= 2992)) || pixel_index == 2998 || pixel_index == 3003 || ((pixel_index >= 3009) && (pixel_index <= 3015)) || pixel_index == 3021 || pixel_index == 3026 || ((pixel_index >= 3034) && (pixel_index <= 3035)) || pixel_index == 3044 || pixel_index == 3049 || ((pixel_index >= 3055) && (pixel_index <= 3056)) || ((pixel_index >= 3060) && (pixel_index <= 3061)) || pixel_index == 3067 || pixel_index == 3076 || ((pixel_index >= 3087) && (pixel_index <= 3088)) || pixel_index == 3094 || pixel_index == 3099 || ((pixel_index >= 3105) && (pixel_index <= 3106)) || pixel_index == 3117 || pixel_index == 3122 || ((pixel_index >= 3130) && (pixel_index <= 3131)) || pixel_index == 3140 || pixel_index == 3145 || ((pixel_index >= 3151) && (pixel_index <= 3152)) || ((pixel_index >= 3156) && (pixel_index <= 3157)) || pixel_index == 3163 || pixel_index == 3172 || ((pixel_index >= 3183) && (pixel_index <= 3184)) || pixel_index == 3190 || pixel_index == 3195 || ((pixel_index >= 3201) && (pixel_index <= 3202)) || pixel_index == 3213 || pixel_index == 3218 || ((pixel_index >= 3226) && (pixel_index <= 3227)) || pixel_index == 3236 || pixel_index == 3241 || ((pixel_index >= 3247) && (pixel_index <= 3248)) || ((pixel_index >= 3252) && (pixel_index <= 3253)) || pixel_index == 3259 || pixel_index == 3268 || ((pixel_index >= 3279) && (pixel_index <= 3280)) || pixel_index == 3286 || pixel_index == 3291 || ((pixel_index >= 3297) && (pixel_index <= 3298)) || pixel_index == 3309 || pixel_index == 3314 || ((pixel_index >= 3322) && (pixel_index <= 3323)) || pixel_index == 3332 || pixel_index == 3337 || ((pixel_index >= 3343) && (pixel_index <= 3344)) || ((pixel_index >= 3348) && (pixel_index <= 3349)) || pixel_index == 3355 || pixel_index == 3364 || ((pixel_index >= 3370) && (pixel_index <= 3376)) || pixel_index == 3382 || pixel_index == 3387 || ((pixel_index >= 3393) && (pixel_index <= 3399)) || pixel_index == 3405 || pixel_index == 3410 || ((pixel_index >= 3418) && (pixel_index <= 3419)) || pixel_index == 3428 || pixel_index == 3433 || ((pixel_index >= 3439) && (pixel_index <= 3445)) || pixel_index == 3451 || pixel_index == 3460 || ((pixel_index >= 3466) && (pixel_index <= 3472)) || pixel_index == 3478 || pixel_index == 3483 || ((pixel_index >= 3489) && (pixel_index <= 3495)) || pixel_index == 3501 || pixel_index == 3506 || ((pixel_index >= 3514) && (pixel_index <= 3515)) || pixel_index == 3524 || pixel_index == 3529 || ((pixel_index >= 3535) && (pixel_index <= 3541)) || pixel_index == 3547 || pixel_index == 3556 || pixel_index == 3574 || pixel_index == 3579 || pixel_index == 3597 || pixel_index == 3602 || pixel_index == 3620 || pixel_index == 3625 || pixel_index == 3643 || pixel_index == 3652 || pixel_index == 3670 || pixel_index == 3675 || pixel_index == 3693 || pixel_index == 3698 || pixel_index == 3716 || pixel_index == 3721 || pixel_index == 3739 || pixel_index == 3748 || pixel_index == 3766 || pixel_index == 3771 || pixel_index == 3789 || pixel_index == 3794 || pixel_index == 3812 || pixel_index == 3817 || pixel_index == 3835 || ((pixel_index >= 3844) && (pixel_index <= 3862)) || ((pixel_index >= 3867) && (pixel_index <= 3885)) || ((pixel_index >= 3890) && (pixel_index <= 3908)) || ((pixel_index >= 3913) && (pixel_index <= 3931)) || pixel_index == 4134 || ((pixel_index >= 4138) && (pixel_index <= 4139)) || ((pixel_index >= 4143) && (pixel_index <= 4144)) || ((pixel_index >= 4148) && (pixel_index <= 4150)) || pixel_index == 4157 || ((pixel_index >= 4161) && (pixel_index <= 4162)) || ((pixel_index >= 4166) && (pixel_index <= 4167)) || ((pixel_index >= 4171) && (pixel_index <= 4173)) || ((pixel_index >= 4181) && (pixel_index <= 4182)) || ((pixel_index >= 4186) && (pixel_index <= 4187)) || ((pixel_index >= 4191) && (pixel_index <= 4193)) || ((pixel_index >= 4205) && (pixel_index <= 4206)) || ((pixel_index >= 4210) && (pixel_index <= 4211)) || ((pixel_index >= 4215) && (pixel_index <= 4217)) || ((pixel_index >= 4229) && (pixel_index <= 4230)) || pixel_index == 4233 || pixel_index == 4236 || pixel_index == 4238 || pixel_index == 4241 || pixel_index == 4243 || ((pixel_index >= 4252) && (pixel_index <= 4253)) || pixel_index == 4256 || pixel_index == 4259 || pixel_index == 4261 || pixel_index == 4264 || pixel_index == 4266 || pixel_index == 4276 || pixel_index == 4279 || pixel_index == 4281 || pixel_index == 4284 || pixel_index == 4286 || pixel_index == 4300 || pixel_index == 4305 || pixel_index == 4308 || pixel_index == 4310 || pixel_index == 4326 || pixel_index == 4331 || pixel_index == 4334 || pixel_index == 4337 || ((pixel_index >= 4340) && (pixel_index <= 4341)) || pixel_index == 4349 || pixel_index == 4352 || pixel_index == 4355 || pixel_index == 4357 || pixel_index == 4360 || ((pixel_index >= 4363) && (pixel_index <= 4364)) || ((pixel_index >= 4373) && (pixel_index <= 4374)) || pixel_index == 4377 || pixel_index == 4380 || ((pixel_index >= 4383) && (pixel_index <= 4384)) || ((pixel_index >= 4396) && (pixel_index <= 4398)) || pixel_index == 4401 || pixel_index == 4404 || ((pixel_index >= 4407) && (pixel_index <= 4408)) || pixel_index == 4422 || pixel_index == 4426 || pixel_index == 4430 || pixel_index == 4433 || pixel_index == 4438 || pixel_index == 4445 || pixel_index == 4448 || pixel_index == 4451 || pixel_index == 4453 || pixel_index == 4456 || pixel_index == 4461 || pixel_index == 4468 || pixel_index == 4471 || pixel_index == 4473 || pixel_index == 4476 || pixel_index == 4481 || pixel_index == 4492 || pixel_index == 4495 || pixel_index == 4497 || pixel_index == 4500 || pixel_index == 4505 || ((pixel_index >= 4517) && (pixel_index <= 4519)) || ((pixel_index >= 4521) && (pixel_index <= 4524)) || ((pixel_index >= 4527) && (pixel_index <= 4528)) || ((pixel_index >= 4531) && (pixel_index <= 4533)) || ((pixel_index >= 4540) && (pixel_index <= 4542)) || ((pixel_index >= 4545) && (pixel_index <= 4546)) || ((pixel_index >= 4550) && (pixel_index <= 4551)) || ((pixel_index >= 4554) && (pixel_index <= 4556)) || ((pixel_index >= 4565) && (pixel_index <= 4566)) || ((pixel_index >= 4570) && (pixel_index <= 4571)) || ((pixel_index >= 4574) && (pixel_index <= 4576)) || ((pixel_index >= 4589) && (pixel_index <= 4590)) || ((pixel_index >= 4594) && (pixel_index <= 4595)) || (pixel_index >= 4598) && (pixel_index <= 4600)) oled_data = 16'b1111111111111111;
    else if (pixel_index == 2213 || pixel_index == 2215 || pixel_index == 2217 || pixel_index == 2219 || pixel_index == 2221 || pixel_index == 2223 || pixel_index == 2225 || pixel_index == 2227 || pixel_index == 2229 || pixel_index == 2405 || pixel_index == 2409 || pixel_index == 2419 || pixel_index == 2421 || pixel_index == 2597 || pixel_index == 2599 || pixel_index == 2601 || pixel_index == 2603 || pixel_index == 2605 || pixel_index == 2609 || pixel_index == 2611 || pixel_index == 2698 || pixel_index == 2705 || pixel_index == 2707 || pixel_index == 2789 || pixel_index == 2791 || ((pixel_index >= 2796) && (pixel_index <= 2797)) || pixel_index == 2802 || pixel_index == 2804 || pixel_index == 2886 || pixel_index == 2888 || pixel_index == 2897 || pixel_index == 2899 || pixel_index == 2981 || pixel_index == 2983 || pixel_index == 2994 || pixel_index == 3080 || pixel_index == 3082 || pixel_index == 3084 || pixel_index == 3086 || pixel_index == 3093 || pixel_index == 3173 || pixel_index == 3175 || pixel_index == 3179 || pixel_index == 3181 || pixel_index == 3272 || pixel_index == 3274 || pixel_index == 3276 || pixel_index == 3278 || pixel_index == 3281 || pixel_index == 3283 || pixel_index == 3365 || pixel_index == 3367 || pixel_index == 3369 || pixel_index == 3378 || pixel_index == 3464 || pixel_index == 3475 || pixel_index == 3557 || pixel_index == 3560 || pixel_index == 3562 || pixel_index == 3564 || pixel_index == 3566 || pixel_index == 3570 || pixel_index == 3572 || pixel_index == 3654 || pixel_index == 3656 || pixel_index == 3658 || pixel_index == 3663 || pixel_index == 3667 || pixel_index == 3669 || pixel_index == 3749 || pixel_index == 3753 || pixel_index == 3755 || pixel_index == 3757 || pixel_index == 3761 || pixel_index == 3764) oled_data = 16'b0010010110101001;
    else if (pixel_index == 2214 || pixel_index == 2216 || pixel_index == 2218 || pixel_index == 2220 || pixel_index == 2222 || pixel_index == 2224 || pixel_index == 2226 || pixel_index == 2228 || pixel_index == 2309 || pixel_index == 2311 || pixel_index == 2313 || pixel_index == 2315 || pixel_index == 2317 || pixel_index == 2319 || pixel_index == 2321 || pixel_index == 2323 || pixel_index == 2325 || pixel_index == 2406 || pixel_index == 2408 || pixel_index == 2418 || pixel_index == 2501 || pixel_index == 2503 || pixel_index == 2513 || pixel_index == 2515 || pixel_index == 2517 || pixel_index == 2598 || pixel_index == 2600 || pixel_index == 2606 || pixel_index == 2612 || pixel_index == 2693 || pixel_index == 2695 || pixel_index == 2697 || pixel_index == 2699 || pixel_index == 2701 || pixel_index == 2708 || pixel_index == 2790 || pixel_index == 2792 || pixel_index == 2795 || pixel_index == 2798 || pixel_index == 2801 || pixel_index == 2805 || pixel_index == 2889 || pixel_index == 2900 || pixel_index == 2982 || pixel_index == 2984 || pixel_index == 2993 || pixel_index == 2995 || pixel_index == 2997 || pixel_index == 3077 || pixel_index == 3079 || pixel_index == 3081 || pixel_index == 3090 || pixel_index == 3092 || pixel_index == 3180 || pixel_index == 3185 || pixel_index == 3187 || pixel_index == 3189 || pixel_index == 3269 || pixel_index == 3271 || pixel_index == 3273 || pixel_index == 3284 || pixel_index == 3366 || pixel_index == 3377 || pixel_index == 3379 || pixel_index == 3381 || pixel_index == 3461 || pixel_index == 3463 || pixel_index == 3465 || pixel_index == 3476 || pixel_index == 3558 || pixel_index == 3563 || pixel_index == 3565 || pixel_index == 3569 || pixel_index == 3655 || pixel_index == 3664 || pixel_index == 3666 || pixel_index == 3668 || pixel_index == 3750 || pixel_index == 3754 || pixel_index == 3756 || pixel_index == 3758 || pixel_index == 3760 || pixel_index == 3762) oled_data = 16'b0010010101101001;
    else if (pixel_index == 2236 || pixel_index == 2238 || pixel_index == 2240 || pixel_index == 2242 || pixel_index == 2246 || pixel_index == 2248 || pixel_index == 2250 || pixel_index == 2252 || pixel_index == 2334 || pixel_index == 2336 || ((pixel_index >= 2340) && (pixel_index <= 2341)) || pixel_index == 2343 || pixel_index == 2345 || pixel_index == 2428 || pixel_index == 2431 || pixel_index == 2441 || pixel_index == 2444 || pixel_index == 2526 || pixel_index == 2528 || pixel_index == 2536 || ((pixel_index >= 2538) && (pixel_index <= 2539)) || pixel_index == 2621 || pixel_index == 2623 || ((pixel_index >= 2625) && (pixel_index <= 2626)) || pixel_index == 2628 || pixel_index == 2633 || pixel_index == 2636 || pixel_index == 2716 || ((pixel_index >= 2719) && (pixel_index <= 2720)) || pixel_index == 2722 || ((pixel_index >= 2724) && (pixel_index <= 2725)) || pixel_index == 2732 || pixel_index == 2813 || ((pixel_index >= 2818) && (pixel_index <= 2819)) || pixel_index == 2821 || pixel_index == 2824 || pixel_index == 2826 || pixel_index == 2910 || pixel_index == 2912 || pixel_index == 2922 || pixel_index == 2924 || pixel_index == 3004 || pixel_index == 3007 || pixel_index == 3016 || pixel_index == 3020 || pixel_index == 3103 || pixel_index == 3107 || pixel_index == 3109 || pixel_index == 3115 || pixel_index == 3196 || pixel_index == 3199 || pixel_index == 3204 || pixel_index == 3206 || ((pixel_index >= 3208) && (pixel_index <= 3209)) || pixel_index == 3212 || pixel_index == 3292 || pixel_index == 3294 || pixel_index == 3300 || pixel_index == 3303 || pixel_index == 3305 || pixel_index == 3308 || pixel_index == 3388 || pixel_index == 3390 || pixel_index == 3392 || pixel_index == 3400 || pixel_index == 3402 || pixel_index == 3487 || ((pixel_index >= 3580) && (pixel_index <= 3581)) || pixel_index == 3583 || pixel_index == 3585 || pixel_index == 3587 || pixel_index == 3589 || pixel_index == 3592 || pixel_index == 3595 || pixel_index == 3677 || pixel_index == 3680 || pixel_index == 3682 || ((pixel_index >= 3685) && (pixel_index <= 3686)) || pixel_index == 3690 || pixel_index == 3772 || ((pixel_index >= 3776) && (pixel_index <= 3777)) || pixel_index == 3779 || pixel_index == 3784 || pixel_index == 3787) oled_data = 16'b1111111000100010;
    else if (pixel_index == 2237 || pixel_index == 2241 || pixel_index == 2243 || pixel_index == 2245 || pixel_index == 2247 || pixel_index == 2251 || pixel_index == 2332 || pixel_index == 2335 || pixel_index == 2338 || pixel_index == 2346 || pixel_index == 2348 || pixel_index == 2429 || pixel_index == 2440 || pixel_index == 2443 || pixel_index == 2525 || pixel_index == 2527 || pixel_index == 2620 || pixel_index == 2627 || pixel_index == 2632 || pixel_index == 2634 || pixel_index == 2718 || pixel_index == 2729 || pixel_index == 2731 || pixel_index == 2812 || pixel_index == 2815 || pixel_index == 2817 || pixel_index == 2825 || pixel_index == 2827 || pixel_index == 2909 || pixel_index == 2911 || pixel_index == 2920 || pixel_index == 3005 || pixel_index == 3017 || pixel_index == 3019 || pixel_index == 3100 || pixel_index == 3102 || pixel_index == 3104 || pixel_index == 3110 || pixel_index == 3112 || pixel_index == 3114 || pixel_index == 3197 || pixel_index == 3203 || pixel_index == 3207 || pixel_index == 3210 || ((pixel_index >= 3295) && (pixel_index <= 3296)) || pixel_index == 3301 || pixel_index == 3307 || pixel_index == 3389 || pixel_index == 3401 || pixel_index == 3403 || pixel_index == 3484 || pixel_index == 3486 || pixel_index == 3496 || pixel_index == 3498 || pixel_index == 3500 || pixel_index == 3584 || pixel_index == 3586 || pixel_index == 3590 || pixel_index == 3593 || pixel_index == 3596 || pixel_index == 3678 || pixel_index == 3684 || pixel_index == 3687 || pixel_index == 3689 || pixel_index == 3691 || pixel_index == 3773 || pixel_index == 3775 || pixel_index == 3778 || pixel_index == 3781 || pixel_index == 3783 || pixel_index == 3786 || pixel_index == 3788) oled_data = 16'b1111110111100010;
    else if (pixel_index == 2239 || pixel_index == 2249 || pixel_index == 2342 || pixel_index == 2432 || pixel_index == 2537 || pixel_index == 2540 || pixel_index == 2622 || pixel_index == 2624 || pixel_index == 2629 || pixel_index == 2721 || pixel_index == 2723 || pixel_index == 2820 || pixel_index == 2923 || pixel_index == 3008 || pixel_index == 3108 || pixel_index == 3116 || pixel_index == 3205 || pixel_index == 3293 || pixel_index == 3304 || pixel_index == 3488 || pixel_index == 3582 || pixel_index == 3588 || pixel_index == 3676 || pixel_index == 3681) oled_data = 16'b1111110111100001;
    else if (pixel_index == 2244 || pixel_index == 2333 || pixel_index == 2337 || pixel_index == 2339 || pixel_index == 2344 || pixel_index == 2347 || pixel_index == 2430 || pixel_index == 2442 || pixel_index == 2524 || pixel_index == 2635 || pixel_index == 2717 || pixel_index == 2728 || pixel_index == 2730 || pixel_index == 2814 || pixel_index == 2816 || pixel_index == 2828 || pixel_index == 2908 || pixel_index == 2921 || pixel_index == 3006 || pixel_index == 3018 || pixel_index == 3101 || pixel_index == 3111 || pixel_index == 3113 || pixel_index == 3198 || pixel_index == 3200 || pixel_index == 3211 || pixel_index == 3299 || pixel_index == 3302 || pixel_index == 3306 || pixel_index == 3391 || pixel_index == 3404 || pixel_index == 3485 || pixel_index == 3497 || pixel_index == 3499 || pixel_index == 3591 || pixel_index == 3594 || pixel_index == 3679 || pixel_index == 3683 || pixel_index == 3688 || pixel_index == 3692 || pixel_index == 3774 || pixel_index == 3780 || pixel_index == 3782 || pixel_index == 3785) oled_data = 16'b1111111000100001;
    else if (((pixel_index >= 2259) && (pixel_index <= 2260)) || ((pixel_index >= 2262) && (pixel_index <= 2264)) || ((pixel_index >= 2266) && (pixel_index <= 2268)) || ((pixel_index >= 2270) && (pixel_index <= 2272)) || ((pixel_index >= 2274) && (pixel_index <= 2275)) || ((pixel_index >= 2356) && (pixel_index <= 2357)) || pixel_index == 2359 || ((pixel_index >= 2361) && (pixel_index <= 2362)) || ((pixel_index >= 2364) && (pixel_index <= 2365)) || pixel_index == 2367 || ((pixel_index >= 2369) && (pixel_index <= 2370)) || ((pixel_index >= 2451) && (pixel_index <= 2452)) || ((pixel_index >= 2454) && (pixel_index <= 2456)) || pixel_index == 2460 || ((pixel_index >= 2462) && (pixel_index <= 2464)) || ((pixel_index >= 2466) && (pixel_index <= 2467)) || pixel_index == 2547 || ((pixel_index >= 2549) && (pixel_index <= 2550)) || ((pixel_index >= 2552) && (pixel_index <= 2553)) || ((pixel_index >= 2556) && (pixel_index <= 2557)) || ((pixel_index >= 2559) && (pixel_index <= 2561)) || pixel_index == 2563 || ((pixel_index >= 2643) && (pixel_index <= 2644)) || ((pixel_index >= 2646) && (pixel_index <= 2647)) || pixel_index == 2649 || ((pixel_index >= 2653) && (pixel_index <= 2654)) || pixel_index == 2656 || ((pixel_index >= 2658) && (pixel_index <= 2659)) || ((pixel_index >= 2740) && (pixel_index <= 2741)) || ((pixel_index >= 2743) && (pixel_index <= 2744)) || ((pixel_index >= 2748) && (pixel_index <= 2749)) || ((pixel_index >= 2751) && (pixel_index <= 2753)) || pixel_index == 2755 || pixel_index == 2835 || ((pixel_index >= 2837) && (pixel_index <= 2838)) || ((pixel_index >= 2840) && (pixel_index <= 2841)) || pixel_index == 2844 || ((pixel_index >= 2846) && (pixel_index <= 2847)) || ((pixel_index >= 2849) && (pixel_index <= 2850)) || ((pixel_index >= 2931) && (pixel_index <= 2932)) || ((pixel_index >= 2934) && (pixel_index <= 2936)) || ((pixel_index >= 2940) && (pixel_index <= 2941)) || ((pixel_index >= 2943) && (pixel_index <= 2944)) || ((pixel_index >= 2946) && (pixel_index <= 2947)) || pixel_index == 3027 || ((pixel_index >= 3029) && (pixel_index <= 3030)) || ((pixel_index >= 3032) && (pixel_index <= 3033)) || ((pixel_index >= 3037) && (pixel_index <= 3038)) || ((pixel_index >= 3040) && (pixel_index <= 3041)) || pixel_index == 3043 || ((pixel_index >= 3123) && (pixel_index <= 3124)) || ((pixel_index >= 3126) && (pixel_index <= 3127)) || pixel_index == 3129 || pixel_index == 3132 || ((pixel_index >= 3134) && (pixel_index <= 3135)) || ((pixel_index >= 3137) && (pixel_index <= 3138)) || ((pixel_index >= 3220) && (pixel_index <= 3221)) || ((pixel_index >= 3223) && (pixel_index <= 3224)) || ((pixel_index >= 3228) && (pixel_index <= 3229)) || ((pixel_index >= 3231) && (pixel_index <= 3232)) || ((pixel_index >= 3234) && (pixel_index <= 3235)) || ((pixel_index >= 3315) && (pixel_index <= 3316)) || ((pixel_index >= 3318) && (pixel_index <= 3319)) || pixel_index == 3321 || pixel_index == 3324 || ((pixel_index >= 3326) && (pixel_index <= 3327)) || ((pixel_index >= 3329) && (pixel_index <= 3330)) || pixel_index == 3411 || ((pixel_index >= 3413) && (pixel_index <= 3414)) || ((pixel_index >= 3416) && (pixel_index <= 3417)) || ((pixel_index >= 3420) && (pixel_index <= 3421)) || ((pixel_index >= 3423) && (pixel_index <= 3425)) || pixel_index == 3427 || ((pixel_index >= 3507) && (pixel_index <= 3508)) || ((pixel_index >= 3510) && (pixel_index <= 3512)) || ((pixel_index >= 3517) && (pixel_index <= 3518)) || pixel_index == 3520 || ((pixel_index >= 3522) && (pixel_index <= 3523)) || ((pixel_index >= 3604) && (pixel_index <= 3605)) || pixel_index == 3607 || ((pixel_index >= 3609) && (pixel_index <= 3612)) || ((pixel_index >= 3614) && (pixel_index <= 3617)) || pixel_index == 3619 || ((pixel_index >= 3699) && (pixel_index <= 3700)) || ((pixel_index >= 3702) && (pixel_index <= 3705)) || pixel_index == 3707 || ((pixel_index >= 3709) && (pixel_index <= 3710)) || pixel_index == 3712 || ((pixel_index >= 3714) && (pixel_index <= 3715)) || pixel_index == 3795 || ((pixel_index >= 3797) && (pixel_index <= 3798)) || pixel_index == 3800 || ((pixel_index >= 3802) && (pixel_index <= 3804)) || ((pixel_index >= 3806) && (pixel_index <= 3807)) || (pixel_index >= 3809) && (pixel_index <= 3810)) oled_data = 16'b1111101111000000;
    else if (pixel_index == 2261 || pixel_index == 2265 || pixel_index == 2269 || pixel_index == 2273 || pixel_index == 2355 || pixel_index == 2358 || pixel_index == 2360 || pixel_index == 2363 || pixel_index == 2366 || pixel_index == 2368 || pixel_index == 2371 || pixel_index == 2453 || pixel_index == 2457 || pixel_index == 2461 || pixel_index == 2465 || pixel_index == 2548 || pixel_index == 2551 || pixel_index == 2558 || pixel_index == 2562 || pixel_index == 2645 || pixel_index == 2648 || pixel_index == 2652 || pixel_index == 2655 || pixel_index == 2657 || pixel_index == 2739 || pixel_index == 2742 || pixel_index == 2745 || pixel_index == 2750 || pixel_index == 2754 || pixel_index == 2836 || pixel_index == 2839 || pixel_index == 2845 || pixel_index == 2848 || pixel_index == 2851 || pixel_index == 2933 || pixel_index == 2937 || pixel_index == 2942 || pixel_index == 2945 || pixel_index == 3028 || pixel_index == 3031 || pixel_index == 3036 || pixel_index == 3039 || pixel_index == 3042 || pixel_index == 3125 || pixel_index == 3128 || pixel_index == 3133 || pixel_index == 3136 || pixel_index == 3139 || pixel_index == 3219 || pixel_index == 3222 || pixel_index == 3225 || pixel_index == 3230 || pixel_index == 3233 || pixel_index == 3317 || pixel_index == 3320 || pixel_index == 3325 || pixel_index == 3328 || pixel_index == 3331 || pixel_index == 3412 || pixel_index == 3415 || pixel_index == 3422 || pixel_index == 3426 || pixel_index == 3509 || pixel_index == 3513 || pixel_index == 3516 || pixel_index == 3519 || pixel_index == 3521 || pixel_index == 3603 || pixel_index == 3606 || pixel_index == 3608 || pixel_index == 3613 || pixel_index == 3618 || pixel_index == 3701 || pixel_index == 3706 || pixel_index == 3708 || pixel_index == 3711 || pixel_index == 3713 || pixel_index == 3796 || pixel_index == 3799 || pixel_index == 3801 || pixel_index == 3805 || pixel_index == 3808 || pixel_index == 3811) oled_data = 16'b1111110000000000;
    else if (pixel_index == 2282 || pixel_index == 2284 || pixel_index == 2287 || pixel_index == 2291 || pixel_index == 2294 || ((pixel_index >= 2296) && (pixel_index <= 2297)) || pixel_index == 2378 || pixel_index == 2381 || pixel_index == 2385 || pixel_index == 2388 || ((pixel_index >= 2390) && (pixel_index <= 2391)) || ((pixel_index >= 2393) && (pixel_index <= 2394)) || pixel_index == 2475 || pixel_index == 2477 || pixel_index == 2488 || pixel_index == 2570 || pixel_index == 2574 || pixel_index == 2582 || pixel_index == 2584 || pixel_index == 2586 || pixel_index == 2667 || pixel_index == 2673 || pixel_index == 2675 || pixel_index == 2680 || pixel_index == 2777 || pixel_index == 2858 || pixel_index == 2860 || ((pixel_index >= 2865) && (pixel_index <= 2867)) || pixel_index == 2870 || pixel_index == 2872 || pixel_index == 2874 || pixel_index == 2958 || pixel_index == 2967 || pixel_index == 3051 || pixel_index == 3057 || pixel_index == 3059 || pixel_index == 3062 || ((pixel_index >= 3064) && (pixel_index <= 3065)) || ((pixel_index >= 3149) && (pixel_index <= 3150)) || pixel_index == 3158 || pixel_index == 3242 || pixel_index == 3249 || pixel_index == 3257 || pixel_index == 3341 || pixel_index == 3347 || pixel_index == 3354 || pixel_index == 3448 || pixel_index == 3530 || pixel_index == 3544 || pixel_index == 3627 || pixel_index == 3633 || pixel_index == 3637 || pixel_index == 3640 || pixel_index == 3722 || pixel_index == 3724 || pixel_index == 3726 || ((pixel_index >= 3729) && (pixel_index <= 3730)) || pixel_index == 3732 || pixel_index == 3734 || pixel_index == 3737 || pixel_index == 3818 || pixel_index == 3821 || pixel_index == 3823 || pixel_index == 3825 || pixel_index == 3827 || pixel_index == 3829 || pixel_index == 3831 || pixel_index == 3833) oled_data = 16'b1110100011000100;
    else if (pixel_index == 2283 || pixel_index == 2295 || pixel_index == 2298 || pixel_index == 2474 || pixel_index == 2476 || pixel_index == 2478 || pixel_index == 2489 || pixel_index == 2585 || pixel_index == 2674 || pixel_index == 2769 || pixel_index == 2771 || pixel_index == 2859 || pixel_index == 2873 || pixel_index == 2961 || pixel_index == 2963 || pixel_index == 3052 || pixel_index == 3054 || pixel_index == 3058 || pixel_index == 3063 || pixel_index == 3345 || pixel_index == 3545 || pixel_index == 3626 || pixel_index == 3634 || pixel_index == 3636 || pixel_index == 3731 || pixel_index == 3738 || pixel_index == 3822 || pixel_index == 3824 || pixel_index == 3830 || pixel_index == 3832) oled_data = 16'b1110100100000101;
    else if (pixel_index == 2285 || pixel_index == 2288 || pixel_index == 2290 || pixel_index == 2293 || pixel_index == 2379 || pixel_index == 2382 || pixel_index == 2384 || pixel_index == 2387 || pixel_index == 2487 || pixel_index == 2572 || pixel_index == 2666 || pixel_index == 2669 || pixel_index == 2678 || pixel_index == 2765 || pixel_index == 2778 || pixel_index == 2862 || pixel_index == 2871 || pixel_index == 2954 || pixel_index == 2956 || pixel_index == 3066 || pixel_index == 3146 || pixel_index == 3148 || pixel_index == 3155 || pixel_index == 3161 || pixel_index == 3243 || pixel_index == 3245 || pixel_index == 3255 || pixel_index == 3258 || pixel_index == 3339 || pixel_index == 3342 || pixel_index == 3346 || pixel_index == 3350 || pixel_index == 3352 || pixel_index == 3434 || pixel_index == 3436 || pixel_index == 3438 || pixel_index == 3447 || pixel_index == 3449 || pixel_index == 3532 || pixel_index == 3542 || pixel_index == 3629 || pixel_index == 3631 || pixel_index == 3639 || pixel_index == 3642 || pixel_index == 3819) oled_data = 16'b1110100100000100;
    else if (pixel_index == 2286 || pixel_index == 2289 || pixel_index == 2292 || pixel_index == 2486 || pixel_index == 2668 || pixel_index == 2670 || pixel_index == 2679 || pixel_index == 2682 || pixel_index == 2762 || pixel_index == 2764 || pixel_index == 2774 || pixel_index == 2776 || pixel_index == 2861 || pixel_index == 2957 || pixel_index == 2968 || pixel_index == 2970 || pixel_index == 3050 || pixel_index == 3154 || pixel_index == 3160 || pixel_index == 3244 || pixel_index == 3250 || pixel_index == 3254 || pixel_index == 3256 || pixel_index == 3338 || pixel_index == 3435 || pixel_index == 3437 || pixel_index == 3446 || pixel_index == 3450 || pixel_index == 3533 || pixel_index == 3628 || pixel_index == 3630 || pixel_index == 3632 || pixel_index == 3638 || pixel_index == 3641 || pixel_index == 3727 || pixel_index == 3735 || pixel_index == 3820 || pixel_index == 3828) oled_data = 16'b1110100011000101;
    else if (pixel_index == 2310 || pixel_index == 2312 || pixel_index == 2314 || pixel_index == 2316 || pixel_index == 2318 || pixel_index == 2320 || pixel_index == 2322 || pixel_index == 2324 || pixel_index == 2502 || pixel_index == 2504 || pixel_index == 2514 || pixel_index == 2516 || pixel_index == 2613 || pixel_index == 2696 || pixel_index == 2700 || pixel_index == 2794 || pixel_index == 2901 || pixel_index == 2985 || pixel_index == 3078 || pixel_index == 3089 || pixel_index == 3091 || pixel_index == 3188 || pixel_index == 3270 || pixel_index == 3380 || pixel_index == 3473 || pixel_index == 3477 || pixel_index == 3559 || pixel_index == 3659 || pixel_index == 3661 || pixel_index == 3665 || pixel_index == 3759) oled_data = 16'b0010010110101010;
    else if (pixel_index == 2380 || pixel_index == 2383 || pixel_index == 2386 || pixel_index == 2571 || pixel_index == 3147 || pixel_index == 3162 || pixel_index == 3246 || pixel_index == 3340 || pixel_index == 3351 || pixel_index == 3353 || pixel_index == 3543) oled_data = 16'b1110000011000101;
    else if (pixel_index == 2389 || pixel_index == 2392 || pixel_index == 2583 || pixel_index == 2966 || pixel_index == 3723 || pixel_index == 3826) oled_data = 16'b1110000100000101;
    else if (pixel_index == 2407 || pixel_index == 2417 || pixel_index == 2709 || pixel_index == 2793 || pixel_index == 2996 || pixel_index == 3177 || pixel_index == 3186 || pixel_index == 3285 || pixel_index == 3568 || pixel_index == 3751) oled_data = 16'b0010110110101001;
    else if (pixel_index == 2420 || pixel_index == 2505 || pixel_index == 2604 || pixel_index == 2610 || pixel_index == 3083 || pixel_index == 3174 || pixel_index == 3182 || pixel_index == 3474 || pixel_index == 3573 || pixel_index == 3657 || pixel_index == 3660 || pixel_index == 3662) oled_data = 16'b0010110101101001;
    else if (pixel_index == 2490 || pixel_index == 2573 || pixel_index == 2766 || pixel_index == 2770 || pixel_index == 2955 || pixel_index == 2962 || pixel_index == 3053 || pixel_index == 3251 || pixel_index == 3531 || pixel_index == 3534 || pixel_index == 3546 || pixel_index == 3635 || pixel_index == 3834) oled_data = 16'b1110000011000100;
    else if (pixel_index == 2602 || pixel_index == 2706 || pixel_index == 2803 || pixel_index == 2885 || pixel_index == 3085 || pixel_index == 3176 || pixel_index == 3178 || pixel_index == 3275 || pixel_index == 3277 || pixel_index == 3282 || pixel_index == 3561 || pixel_index == 3567 || pixel_index == 3571 || pixel_index == 3653 || pixel_index == 3752 || pixel_index == 3765) oled_data = 16'b0010010101101010;
    else if (pixel_index == 2681 || pixel_index == 2763 || pixel_index == 2775 || pixel_index == 2969 || pixel_index == 3153 || pixel_index == 3159 || pixel_index == 3725 || pixel_index == 3728 || pixel_index == 3733 || pixel_index == 3736) oled_data = 16'b1110000100000100;
    else if (pixel_index == 2694 || pixel_index == 2702 || pixel_index == 3462 || pixel_index == 3763) oled_data = 16'b0010110110101010;
    else if (pixel_index == 2887 || pixel_index == 2898 || pixel_index == 3368) oled_data = 16'b0010110101101010;
    else if (pixel_index == 5206 || pixel_index == 5305 || pixel_index == 5307 || pixel_index == 5319 || pixel_index == 5327 || pixel_index == 5341 || pixel_index == 5396 || pixel_index == 5421 || pixel_index == 5430 || pixel_index == 5501 || pixel_index == 5507 || pixel_index == 5606 || pixel_index == 5619 || pixel_index == 5622 || pixel_index == 5634 || pixel_index == 5642 || pixel_index == 5693 || pixel_index == 5695 || pixel_index == 5698 || pixel_index == 5710 || pixel_index == 5732 || pixel_index == 5741) oled_data = 16'b0101001101011110;
    else if (pixel_index == 5260 || pixel_index == 5301 || pixel_index == 5309 || pixel_index == 5314 || pixel_index == 5316 || pixel_index == 5330 || pixel_index == 5336 || pixel_index == 5338 || pixel_index == 5343 || pixel_index == 5347 || pixel_index == 5351 || pixel_index == 5354 || pixel_index == 5417 || pixel_index == 5442 || pixel_index == 5497 || pixel_index == 5511 || pixel_index == 5522 || pixel_index == 5543 || pixel_index == 5545 || pixel_index == 5592 || pixel_index == 5621 || pixel_index == 5625 || pixel_index == 5630 || pixel_index == 5646 || pixel_index == 5714 || pixel_index == 5782 || pixel_index == 5836) oled_data = 16'b0100101101011110;
    else if (pixel_index == 5304 || pixel_index == 5306 || pixel_index == 5318 || pixel_index == 5320 || pixel_index == 5326 || pixel_index == 5328 || pixel_index == 5334 || pixel_index == 5340 || pixel_index == 5342 || pixel_index == 5357 || pixel_index == 5492 || pixel_index == 5510 || pixel_index == 5518 || pixel_index == 5524 || pixel_index == 5550 || pixel_index == 5597 || pixel_index == 5603 || pixel_index == 5618 || pixel_index == 5637 || pixel_index == 5696 || pixel_index == 5709 || pixel_index == 5720 || pixel_index == 5722 || pixel_index == 5731 || pixel_index == 5738) oled_data = 16'b0100101101011101;
    else if (pixel_index == 5315 || pixel_index == 5337 || pixel_index == 5344 || pixel_index == 5348 || pixel_index == 5447 || pixel_index == 5450 || pixel_index == 5496 || pixel_index == 5529 || pixel_index == 5534 || pixel_index == 5616 || pixel_index == 5639 || pixel_index == 5685 || pixel_index == 5700) oled_data = 16'b0101001101011101;
    else if (pixel_index == 5400 || pixel_index == 5433 || pixel_index == 5438 || pixel_index == 5445 || pixel_index == 5519 || pixel_index == 5588 || pixel_index == 5699 || pixel_index == 5735) oled_data = 16'b0100101110011110;
    else if (pixel_index == 5405 || pixel_index == 5411 || pixel_index == 5498 || pixel_index == 5526 || pixel_index == 5538 || pixel_index == 5544 || pixel_index == 5546 || pixel_index == 5688 || pixel_index == 5694 || pixel_index == 5702 || pixel_index == 5711 || pixel_index == 5718 || pixel_index == 5726) oled_data = 16'b0100101110011101;
    else if (pixel_index == 5414 || pixel_index == 5454 || pixel_index == 5721) oled_data = 16'b0101001110011110;
    else if (pixel_index == 5426 || pixel_index == 5512) oled_data = 16'b0101001110011101;
    else oled_data = 0;




    end

endmodule