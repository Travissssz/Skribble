`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.04.2025 02:55:51
// Design Name: 
// Module Name: bunny_frame
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bunny_frame(input frame_rate, input [12:0] pixel_index, output reg [15:0] oled_data);
    reg [15:0] frame_count = 1;
    parameter picture_total_count = 1;
    
    always @ (posedge frame_rate) begin
        frame_count <= (frame_count == picture_total_count - 1) ? 0 : frame_count + 1;
    end
   
    always @ (*) begin
        if (((pixel_index >= 0) && (pixel_index <= 96)) || pixel_index == 98 || pixel_index == 100 || pixel_index == 102 || pixel_index == 104 || pixel_index == 106 || pixel_index == 108 || pixel_index == 110 || pixel_index == 112 || pixel_index == 114 || pixel_index == 116 || pixel_index == 118 || pixel_index == 120 || pixel_index == 122 || pixel_index == 124 || pixel_index == 126 || pixel_index == 128 || pixel_index == 130 || pixel_index == 132 || pixel_index == 134 || pixel_index == 136 || pixel_index == 138 || pixel_index == 140 || pixel_index == 142 || pixel_index == 144 || pixel_index == 146 || pixel_index == 148 || pixel_index == 150 || pixel_index == 152 || pixel_index == 154 || pixel_index == 156 || pixel_index == 158 || pixel_index == 160 || pixel_index == 162 || pixel_index == 164 || pixel_index == 166 || pixel_index == 168 || pixel_index == 170 || pixel_index == 172 || pixel_index == 174 || pixel_index == 176 || pixel_index == 178 || pixel_index == 180 || pixel_index == 182 || pixel_index == 184 || pixel_index == 186 || pixel_index == 188 || pixel_index == 190 || ((pixel_index >= 192) && (pixel_index <= 195)) || ((pixel_index >= 197) && (pixel_index <= 201)) || ((pixel_index >= 203) && (pixel_index <= 207)) || ((pixel_index >= 209) && (pixel_index <= 213)) || ((pixel_index >= 215) && (pixel_index <= 219)) || ((pixel_index >= 221) && (pixel_index <= 225)) || ((pixel_index >= 227) && (pixel_index <= 231)) || ((pixel_index >= 233) && (pixel_index <= 237)) || ((pixel_index >= 239) && (pixel_index <= 240)) || ((pixel_index >= 248) && (pixel_index <= 251)) || ((pixel_index >= 253) && (pixel_index <= 257)) || ((pixel_index >= 259) && (pixel_index <= 263)) || ((pixel_index >= 265) && (pixel_index <= 269)) || ((pixel_index >= 271) && (pixel_index <= 275)) || ((pixel_index >= 277) && (pixel_index <= 281)) || ((pixel_index >= 283) && (pixel_index <= 286)) || pixel_index == 288 || pixel_index == 292 || pixel_index == 298 || pixel_index == 304 || pixel_index == 310 || pixel_index == 316 || pixel_index == 334 || pixel_index == 346 || pixel_index == 348 || pixel_index == 354 || pixel_index == 360 || pixel_index == 366 || pixel_index == 372 || pixel_index == 378 || ((pixel_index >= 384) && (pixel_index <= 392)) || ((pixel_index >= 394) && (pixel_index <= 398)) || ((pixel_index >= 400) && (pixel_index <= 404)) || ((pixel_index >= 406) && (pixel_index <= 410)) || ((pixel_index >= 412) && (pixel_index <= 416)) || ((pixel_index >= 426) && (pixel_index <= 428)) || pixel_index == 430 || ((pixel_index >= 442) && (pixel_index <= 448)) || ((pixel_index >= 450) && (pixel_index <= 454)) || ((pixel_index >= 456) && (pixel_index <= 460)) || ((pixel_index >= 462) && (pixel_index <= 466)) || ((pixel_index >= 468) && (pixel_index <= 472)) || ((pixel_index >= 474) && (pixel_index <= 477)) || pixel_index == 480 || pixel_index == 482 || pixel_index == 484 || pixel_index == 486 || pixel_index == 488 || pixel_index == 496 || pixel_index == 498 || pixel_index == 500 || pixel_index == 508 || pixel_index == 510 || pixel_index == 524 || pixel_index == 526 || pixel_index == 573 || ((pixel_index >= 575) && (pixel_index <= 583)) || ((pixel_index >= 585) && (pixel_index <= 591)) || ((pixel_index >= 593) && (pixel_index <= 595)) || ((pixel_index >= 597) && (pixel_index <= 603)) || ((pixel_index >= 605) && (pixel_index <= 606)) || ((pixel_index >= 619) && (pixel_index <= 620)) || ((pixel_index >= 635) && (pixel_index <= 638)) || ((pixel_index >= 640) && (pixel_index <= 647)) || ((pixel_index >= 649) && (pixel_index <= 651)) || ((pixel_index >= 653) && (pixel_index <= 659)) || ((pixel_index >= 661) && (pixel_index <= 663)) || ((pixel_index >= 665) && (pixel_index <= 668)) || pixel_index == 670 || pixel_index == 672 || pixel_index == 674 || pixel_index == 678 || pixel_index == 680 || pixel_index == 692 || pixel_index == 718 || pixel_index == 732 || pixel_index == 734 || pixel_index == 744 || pixel_index == 756 || pixel_index == 764 || pixel_index == 766 || ((pixel_index >= 768) && (pixel_index <= 771)) || ((pixel_index >= 773) && (pixel_index <= 774)) || pixel_index == 776 || ((pixel_index >= 778) && (pixel_index <= 783)) || ((pixel_index >= 785) && (pixel_index <= 787)) || ((pixel_index >= 789) && (pixel_index <= 795)) || pixel_index == 797 || pixel_index == 813 || ((pixel_index >= 828) && (pixel_index <= 829)) || ((pixel_index >= 831) && (pixel_index <= 838)) || ((pixel_index >= 840) && (pixel_index <= 843)) || ((pixel_index >= 845) && (pixel_index <= 851)) || ((pixel_index >= 853) && (pixel_index <= 855)) || ((pixel_index >= 857) && (pixel_index <= 858)) || pixel_index == 860 || pixel_index == 862 || pixel_index == 864 || pixel_index == 866 || pixel_index == 868 || pixel_index == 870 || pixel_index == 872 || pixel_index == 874 || pixel_index == 876 || pixel_index == 878 || pixel_index == 880 || pixel_index == 882 || pixel_index == 884 || ((pixel_index >= 892) && (pixel_index <= 893)) || pixel_index == 908 || pixel_index == 910 || pixel_index == 924 || pixel_index == 926 || pixel_index == 934 || pixel_index == 940 || pixel_index == 948 || pixel_index == 952 || pixel_index == 954 || pixel_index == 956 || pixel_index == 958 || ((pixel_index >= 960) && (pixel_index <= 964)) || pixel_index == 966 || pixel_index == 968 || ((pixel_index >= 970) && (pixel_index <= 973)) || ((pixel_index >= 975) && (pixel_index <= 977)) || pixel_index == 979 || ((pixel_index >= 981) && (pixel_index <= 986)) || pixel_index == 1004 || pixel_index == 1006 || pixel_index == 1021 || ((pixel_index >= 1023) && (pixel_index <= 1028)) || ((pixel_index >= 1030) && (pixel_index <= 1034)) || ((pixel_index >= 1036) && (pixel_index <= 1042)) || ((pixel_index >= 1044) && (pixel_index <= 1046)) || pixel_index == 1048 || pixel_index == 1050 || pixel_index == 1052 || pixel_index == 1056 || pixel_index == 1060 || pixel_index == 1062 || pixel_index == 1072 || pixel_index == 1074 || pixel_index == 1078 || pixel_index == 1080 || ((pixel_index >= 1084) && (pixel_index <= 1085)) || pixel_index == 1101 || pixel_index == 1116 || pixel_index == 1118 || pixel_index == 1122 || pixel_index == 1124 || pixel_index == 1130 || pixel_index == 1142 || pixel_index == 1146 || pixel_index == 1148 || pixel_index == 1150 || ((pixel_index >= 1152) && (pixel_index <= 1155)) || pixel_index == 1157 || ((pixel_index >= 1161) && (pixel_index <= 1167)) || pixel_index == 1169 || ((pixel_index >= 1171) && (pixel_index <= 1177)) || pixel_index == 1179 || pixel_index == 1197 || pixel_index == 1212 || pixel_index == 1214 || ((pixel_index >= 1216) && (pixel_index <= 1219)) || ((pixel_index >= 1221) && (pixel_index <= 1224)) || ((pixel_index >= 1226) && (pixel_index <= 1232)) || ((pixel_index >= 1234) && (pixel_index <= 1236)) || pixel_index == 1238 || pixel_index == 1240 || pixel_index == 1242 || pixel_index == 1244 || pixel_index == 1246 || pixel_index == 1248 || pixel_index == 1250 || pixel_index == 1252 || pixel_index == 1254 || pixel_index == 1256 || ((pixel_index >= 1276) && (pixel_index <= 1277)) || ((pixel_index >= 1293) && (pixel_index <= 1294)) || pixel_index == 1308 || pixel_index == 1310 || pixel_index == 1312 || pixel_index == 1314 || pixel_index == 1316 || pixel_index == 1320 || pixel_index == 1330 || pixel_index == 1332 || pixel_index == 1334 || pixel_index == 1336 || pixel_index == 1338 || pixel_index == 1340 || pixel_index == 1342 || ((pixel_index >= 1344) && (pixel_index <= 1348)) || pixel_index == 1350 || ((pixel_index >= 1353) && (pixel_index <= 1360)) || ((pixel_index >= 1362) && (pixel_index <= 1367)) || pixel_index == 1369 || pixel_index == 1371 || pixel_index == 1404 || ((pixel_index >= 1406) && (pixel_index <= 1409)) || pixel_index == 1411 || ((pixel_index >= 1413) && (pixel_index <= 1414)) || pixel_index == 1416 || ((pixel_index >= 1418) && (pixel_index <= 1425)) || ((pixel_index >= 1427) && (pixel_index <= 1428)) || pixel_index == 1430 || pixel_index == 1432 || pixel_index == 1434 || pixel_index == 1436 || pixel_index == 1438 || pixel_index == 1440 || pixel_index == 1442 || pixel_index == 1448 || pixel_index == 1452 || pixel_index == 1454 || pixel_index == 1458 || pixel_index == 1460 || pixel_index == 1464 || pixel_index == 1466 || pixel_index == 1468 || pixel_index == 1470 || ((pixel_index >= 1485) && (pixel_index <= 1486)) || pixel_index == 1507 || pixel_index == 1513 || pixel_index == 1525 || pixel_index == 1527 || pixel_index == 1531 || pixel_index == 1533 || ((pixel_index >= 1535) && (pixel_index <= 1539)) || pixel_index == 1541 || ((pixel_index >= 1543) && (pixel_index <= 1550)) || ((pixel_index >= 1553) && (pixel_index <= 1556)) || ((pixel_index >= 1558) && (pixel_index <= 1560)) || pixel_index == 1562 || pixel_index == 1564 || pixel_index == 1566 || ((pixel_index >= 1597) && (pixel_index <= 1601)) || ((pixel_index >= 1603) && (pixel_index <= 1606)) || pixel_index == 1608 || ((pixel_index >= 1610) && (pixel_index <= 1614)) || ((pixel_index >= 1616) && (pixel_index <= 1618)) || pixel_index == 1620 || pixel_index == 1622 || pixel_index == 1624 || pixel_index == 1626 || ((pixel_index >= 1631) && (pixel_index <= 1632)) || pixel_index == 1634 || pixel_index == 1636 || pixel_index == 1646 || pixel_index == 1648 || pixel_index == 1650 || pixel_index == 1652 || pixel_index == 1654 || pixel_index == 1656 || pixel_index == 1658 || pixel_index == 1660 || pixel_index == 1662 || pixel_index == 1692 || pixel_index == 1704 || pixel_index == 1706 || pixel_index == 1708 || pixel_index == 1710 || pixel_index == 1712 || pixel_index == 1714 || pixel_index == 1716 || pixel_index == 1718 || pixel_index == 1720 || pixel_index == 1722 || pixel_index == 1724 || pixel_index == 1726 || ((pixel_index >= 1728) && (pixel_index <= 1729)) || pixel_index == 1731 || ((pixel_index >= 1733) && (pixel_index <= 1741)) || ((pixel_index >= 1743) && (pixel_index <= 1751)) || pixel_index == 1753 || pixel_index == 1755 || pixel_index == 1757 || pixel_index == 1774 || pixel_index == 1788 || pixel_index == 1790 || ((pixel_index >= 1792) && (pixel_index <= 1793)) || ((pixel_index >= 1795) && (pixel_index <= 1797)) || pixel_index == 1799 || pixel_index == 1801 || ((pixel_index >= 1803) && (pixel_index <= 1809)) || pixel_index == 1811 || pixel_index == 1813 || pixel_index == 1815 || pixel_index == 1817 || pixel_index == 1821 || ((pixel_index >= 1823) && (pixel_index <= 1824)) || pixel_index == 1832 || pixel_index == 1834 || pixel_index == 1838 || ((pixel_index >= 1851) && (pixel_index <= 1853)) || pixel_index == 1855 || pixel_index == 1884 || pixel_index == 1886 || pixel_index == 1888 || pixel_index == 1890 || pixel_index == 1896 || pixel_index == 1908 || pixel_index == 1910 || pixel_index == 1912 || pixel_index == 1914 || pixel_index == 1916 || pixel_index == 1918 || ((pixel_index >= 1920) && (pixel_index <= 1922)) || ((pixel_index >= 1924) && (pixel_index <= 1929)) || ((pixel_index >= 1932) && (pixel_index <= 1934)) || ((pixel_index >= 1936) && (pixel_index <= 1940)) || pixel_index == 1942 || pixel_index == 1945 || pixel_index == 1947 || pixel_index == 1949 || ((pixel_index >= 1981) && (pixel_index <= 1983)) || pixel_index == 1985 || ((pixel_index >= 1987) && (pixel_index <= 1989)) || pixel_index == 1991 || pixel_index == 1993 || ((pixel_index >= 1995) && (pixel_index <= 2000)) || pixel_index == 2002 || pixel_index == 2004 || ((pixel_index >= 2006) && (pixel_index <= 2008)) || pixel_index == 2010 || pixel_index == 2012 || pixel_index == 2014 || pixel_index == 2016 || pixel_index == 2018 || pixel_index == 2020 || pixel_index == 2026 || pixel_index == 2030 || pixel_index == 2032 || pixel_index == 2034 || pixel_index == 2036 || pixel_index == 2038 || pixel_index == 2040 || pixel_index == 2042 || pixel_index == 2044 || pixel_index == 2046 || pixel_index == 2079 || pixel_index == 2081 || pixel_index == 2085 || pixel_index == 2087 || pixel_index == 2089 || pixel_index == 2097 || pixel_index == 2103 || pixel_index == 2105 || pixel_index == 2107 || ((pixel_index >= 2111) && (pixel_index <= 2113)) || ((pixel_index >= 2115) && (pixel_index <= 2121)) || ((pixel_index >= 2123) && (pixel_index <= 2124)) || pixel_index == 2126 || ((pixel_index >= 2128) && (pixel_index <= 2131)) || pixel_index == 2140 || pixel_index == 2172 || pixel_index == 2175 || ((pixel_index >= 2177) && (pixel_index <= 2179)) || pixel_index == 2181 || pixel_index == 2183 || ((pixel_index >= 2186) && (pixel_index <= 2190)) || pixel_index == 2195 || ((pixel_index >= 2197) && (pixel_index <= 2199)) || pixel_index == 2201 || ((pixel_index >= 2205) && (pixel_index <= 2208)) || pixel_index == 2210 || pixel_index == 2218 || pixel_index == 2222 || pixel_index == 2228 || pixel_index == 2230 || pixel_index == 2232 || pixel_index == 2234 || pixel_index == 2236 || pixel_index == 2271 || pixel_index == 2277 || pixel_index == 2279 || pixel_index == 2287 || pixel_index == 2289 || pixel_index == 2291 || pixel_index == 2293 || pixel_index == 2295 || pixel_index == 2299 || pixel_index == 2304 || ((pixel_index >= 2306) && (pixel_index <= 2313)) || pixel_index == 2315 || pixel_index == 2317 || ((pixel_index >= 2319) && (pixel_index <= 2323)) || pixel_index == 2325 || pixel_index == 2327 || pixel_index == 2369 || pixel_index == 2371 || pixel_index == 2373 || pixel_index == 2375 || ((pixel_index >= 2377) && (pixel_index <= 2381)) || pixel_index == 2383 || pixel_index == 2387 || pixel_index == 2390 || pixel_index == 2394 || ((pixel_index >= 2397) && (pixel_index <= 2398)) || pixel_index == 2400 || pixel_index == 2412 || pixel_index == 2414 || pixel_index == 2420 || pixel_index == 2422 || pixel_index == 2424 || pixel_index == 2426 || pixel_index == 2463 || pixel_index == 2465 || pixel_index == 2467 || pixel_index == 2469 || pixel_index == 2471 || pixel_index == 2473 || pixel_index == 2475 || pixel_index == 2477 || pixel_index == 2479 || pixel_index == 2481 || pixel_index == 2488 || pixel_index == 2490 || ((pixel_index >= 2495) && (pixel_index <= 2496)) || ((pixel_index >= 2498) && (pixel_index <= 2504)) || pixel_index == 2506 || pixel_index == 2509 || ((pixel_index >= 2511) && (pixel_index <= 2514)) || pixel_index == 2516 || pixel_index == 2561 || pixel_index == 2563 || pixel_index == 2565 || pixel_index == 2567 || ((pixel_index >= 2569) && (pixel_index <= 2572)) || pixel_index == 2574 || pixel_index == 2578 || ((pixel_index >= 2580) && (pixel_index <= 2582)) || pixel_index == 2584 || pixel_index == 2586 || ((pixel_index >= 2588) && (pixel_index <= 2589)) || ((pixel_index >= 2591) && (pixel_index <= 2592)) || pixel_index == 2596 || pixel_index == 2598 || pixel_index == 2600 || pixel_index == 2602 || pixel_index == 2604 || pixel_index == 2608 || pixel_index == 2610 || pixel_index == 2612 || pixel_index == 2614 || pixel_index == 2616 || pixel_index == 2658 || pixel_index == 2660 || pixel_index == 2664 || pixel_index == 2666 || pixel_index == 2668 || pixel_index == 2672 || pixel_index == 2680 || ((pixel_index >= 2687) && (pixel_index <= 2688)) || ((pixel_index >= 2690) && (pixel_index <= 2695)) || pixel_index == 2697 || pixel_index == 2699 || ((pixel_index >= 2701) && (pixel_index <= 2706)) || pixel_index == 2708 || pixel_index == 2710 || pixel_index == 2753 || pixel_index == 2755 || pixel_index == 2757 || pixel_index == 2759 || ((pixel_index >= 2762) && (pixel_index <= 2764)) || pixel_index == 2766 || ((pixel_index >= 2770) && (pixel_index <= 2772)) || pixel_index == 2774 || ((pixel_index >= 2777) && (pixel_index <= 2778)) || pixel_index == 2781 || pixel_index == 2784 || pixel_index == 2786 || pixel_index == 2788 || pixel_index == 2790 || pixel_index == 2794 || pixel_index == 2796 || pixel_index == 2798 || pixel_index == 2800 || pixel_index == 2802 || pixel_index == 2804 || pixel_index == 2856 || pixel_index == 2860 || pixel_index == 2862 || pixel_index == 2864 || pixel_index == 2868 || pixel_index == 2875 || pixel_index == 2877 || ((pixel_index >= 2879) && (pixel_index <= 2880)) || ((pixel_index >= 2882) && (pixel_index <= 2885)) || pixel_index == 2887 || pixel_index == 2889 || pixel_index == 2891 || ((pixel_index >= 2894) && (pixel_index <= 2897)) || pixel_index == 2899 || pixel_index == 2901 || pixel_index == 2903 || pixel_index == 2946 || pixel_index == 2948 || pixel_index == 2950 || ((pixel_index >= 2953) && (pixel_index <= 2954)) || pixel_index == 2956 || pixel_index == 2958 || pixel_index == 2960 || ((pixel_index >= 2962) && (pixel_index <= 2963)) || pixel_index == 2965 || pixel_index == 2967 || pixel_index == 2969 || pixel_index == 2971 || ((pixel_index >= 2975) && (pixel_index <= 2976)) || pixel_index == 2988 || pixel_index == 2996 || pixel_index == 2998 || pixel_index == 3045 || pixel_index == 3047 || pixel_index == 3051 || pixel_index == 3055 || pixel_index == 3057 || pixel_index == 3061 || pixel_index == 3066 || ((pixel_index >= 3068) && (pixel_index <= 3070)) || pixel_index == 3072 || ((pixel_index >= 3074) && (pixel_index <= 3077)) || pixel_index == 3079 || pixel_index == 3081 || pixel_index == 3083 || ((pixel_index >= 3085) && (pixel_index <= 3089)) || pixel_index == 3091 || pixel_index == 3093 || pixel_index == 3095 || pixel_index == 3139 || ((pixel_index >= 3141) && (pixel_index <= 3143)) || ((pixel_index >= 3145) && (pixel_index <= 3146)) || pixel_index == 3148 || pixel_index == 3150 || pixel_index == 3154 || pixel_index == 3156 || ((pixel_index >= 3158) && (pixel_index <= 3160)) || pixel_index == 3163 || ((pixel_index >= 3167) && (pixel_index <= 3168)) || pixel_index == 3170 || pixel_index == 3172 || pixel_index == 3176 || pixel_index == 3178 || pixel_index == 3180 || pixel_index == 3188 || pixel_index == 3234 || pixel_index == 3236 || pixel_index == 3238 || pixel_index == 3240 || pixel_index == 3248 || pixel_index == 3252 || pixel_index == 3257 || ((pixel_index >= 3260) && (pixel_index <= 3261)) || ((pixel_index >= 3263) && (pixel_index <= 3264)) || ((pixel_index >= 3266) && (pixel_index <= 3267)) || pixel_index == 3271 || pixel_index == 3273 || ((pixel_index >= 3277) && (pixel_index <= 3279)) || pixel_index == 3281 || pixel_index == 3283 || ((pixel_index >= 3285) && (pixel_index <= 3287)) || pixel_index == 3330 || ((pixel_index >= 3332) && (pixel_index <= 3334)) || ((pixel_index >= 3336) && (pixel_index <= 3339)) || pixel_index == 3341 || pixel_index == 3343 || pixel_index == 3345 || pixel_index == 3348 || ((pixel_index >= 3350) && (pixel_index <= 3351)) || pixel_index == 3353 || pixel_index == 3357 || pixel_index == 3360 || pixel_index == 3364 || pixel_index == 3366 || pixel_index == 3368 || pixel_index == 3370 || pixel_index == 3372 || pixel_index == 3378 || pixel_index == 3380 || pixel_index == 3382 || pixel_index == 3427 || pixel_index == 3431 || pixel_index == 3435 || pixel_index == 3437 || pixel_index == 3439 || pixel_index == 3443 || pixel_index == 3448 || ((pixel_index >= 3451) && (pixel_index <= 3452)) || ((pixel_index >= 3454) && (pixel_index <= 3456)) || pixel_index == 3458 || pixel_index == 3462 || ((pixel_index >= 3464) && (pixel_index <= 3466)) || ((pixel_index >= 3468) && (pixel_index <= 3471)) || pixel_index == 3473 || pixel_index == 3475 || ((pixel_index >= 3477) && (pixel_index <= 3478)) || pixel_index == 3522 || ((pixel_index >= 3524) && (pixel_index <= 3525)) || ((pixel_index >= 3528) && (pixel_index <= 3530)) || pixel_index == 3532 || ((pixel_index >= 3537) && (pixel_index <= 3538)) || pixel_index == 3540 || pixel_index == 3542 || pixel_index == 3546 || pixel_index == 3548 || pixel_index == 3552 || pixel_index == 3554 || pixel_index == 3556 || pixel_index == 3560 || pixel_index == 3562 || pixel_index == 3618 || pixel_index == 3622 || pixel_index == 3630 || pixel_index == 3634 || pixel_index == 3639 || pixel_index == 3641 || pixel_index == 3643 || ((pixel_index >= 3645) && (pixel_index <= 3646)) || pixel_index == 3648 || pixel_index == 3650 || pixel_index == 3652 || ((pixel_index >= 3654) && (pixel_index <= 3659)) || ((pixel_index >= 3661) && (pixel_index <= 3662)) || pixel_index == 3664 || pixel_index == 3666 || ((pixel_index >= 3668) && (pixel_index <= 3669)) || pixel_index == 3671 || ((pixel_index >= 3715) && (pixel_index <= 3717)) || pixel_index == 3719 || pixel_index == 3722 || pixel_index == 3724 || ((pixel_index >= 3727) && (pixel_index <= 3728)) || pixel_index == 3730 || ((pixel_index >= 3732) && (pixel_index <= 3733)) || pixel_index == 3735 || pixel_index == 3737 || pixel_index == 3739 || pixel_index == 3741 || ((pixel_index >= 3743) && (pixel_index <= 3744)) || pixel_index == 3746 || pixel_index == 3748 || pixel_index == 3750 || pixel_index == 3752 || pixel_index == 3754 || pixel_index == 3756 || pixel_index == 3760 || pixel_index == 3762 || pixel_index == 3767 || pixel_index == 3810 || pixel_index == 3816 || pixel_index == 3820 || pixel_index == 3824 || pixel_index == 3831 || pixel_index == 3833 || pixel_index == 3836 || pixel_index == 3838 || pixel_index == 3840 || pixel_index == 3842 || pixel_index == 3844 || ((pixel_index >= 3846) && (pixel_index <= 3850)) || ((pixel_index >= 3852) && (pixel_index <= 3853)) || pixel_index == 3855 || pixel_index == 3857 || ((pixel_index >= 3860) && (pixel_index <= 3861)) || pixel_index == 3905 || pixel_index == 3908 || pixel_index == 3911 || pixel_index == 3913 || pixel_index == 3915 || pixel_index == 3917 || pixel_index == 3921 || pixel_index == 3923 || pixel_index == 3925 || pixel_index == 3927 || pixel_index == 3929 || pixel_index == 3936 || pixel_index == 3940 || pixel_index == 3950 || pixel_index == 3952 || pixel_index == 3954 || pixel_index == 3956 || ((pixel_index >= 3958) && (pixel_index <= 3959)) || pixel_index == 4000 || pixel_index == 4002 || pixel_index == 4005 || pixel_index == 4007 || pixel_index == 4009 || pixel_index == 4011 || pixel_index == 4015 || pixel_index == 4017 || pixel_index == 4019 || pixel_index == 4021 || pixel_index == 4023 || pixel_index == 4025 || ((pixel_index >= 4027) && (pixel_index <= 4028)) || pixel_index == 4030 || pixel_index == 4032 || ((pixel_index >= 4034) && (pixel_index <= 4035)) || ((pixel_index >= 4037) && (pixel_index <= 4042)) || pixel_index == 4044 || pixel_index == 4046 || pixel_index == 4048 || ((pixel_index >= 4050) && (pixel_index <= 4051)) || pixel_index == 4053 || pixel_index == 4056 || pixel_index == 4097 || pixel_index == 4100 || pixel_index == 4104 || pixel_index == 4106 || ((pixel_index >= 4109) && (pixel_index <= 4110)) || ((pixel_index >= 4112) && (pixel_index <= 4113)) || pixel_index == 4116 || pixel_index == 4118 || pixel_index == 4120 || pixel_index == 4122 || pixel_index == 4126 || pixel_index == 4128 || pixel_index == 4132 || pixel_index == 4144 || pixel_index == 4146 || pixel_index == 4148 || pixel_index == 4150 || pixel_index == 4192 || ((pixel_index >= 4194) && (pixel_index <= 4195)) || pixel_index == 4197 || pixel_index == 4199 || pixel_index == 4201 || pixel_index == 4203 || pixel_index == 4210 || pixel_index == 4212 || ((pixel_index >= 4214) && (pixel_index <= 4215)) || pixel_index == 4219 || pixel_index == 4224 || pixel_index == 4226 || ((pixel_index >= 4229) && (pixel_index <= 4233)) || pixel_index == 4235 || pixel_index == 4237 || pixel_index == 4239 || ((pixel_index >= 4241) && (pixel_index <= 4242)) || ((pixel_index >= 4244) && (pixel_index <= 4245)) || pixel_index == 4247 || pixel_index == 4289 || pixel_index == 4293 || pixel_index == 4295 || pixel_index == 4297 || pixel_index == 4299 || pixel_index == 4301 || pixel_index == 4303 || pixel_index == 4310 || pixel_index == 4312 || pixel_index == 4316 || ((pixel_index >= 4318) && (pixel_index <= 4320)) || pixel_index == 4322 || pixel_index == 4334 || pixel_index == 4336 || pixel_index == 4338 || pixel_index == 4340 || pixel_index == 4342 || ((pixel_index >= 4386) && (pixel_index <= 4387)) || pixel_index == 4400 || pixel_index == 4402 || ((pixel_index >= 4405) && (pixel_index <= 4409)) || pixel_index == 4412 || pixel_index == 4416 || pixel_index == 4418 || pixel_index == 4420 || ((pixel_index >= 4422) && (pixel_index <= 4424)) || ((pixel_index >= 4426) && (pixel_index <= 4427)) || pixel_index == 4430 || ((pixel_index >= 4432) && (pixel_index <= 4434)) || ((pixel_index >= 4437) && (pixel_index <= 4439)) || pixel_index == 4482 || pixel_index == 4484 || pixel_index == 4486 || pixel_index == 4488 || pixel_index == 4490 || ((pixel_index >= 4492) && (pixel_index <= 4493)) || pixel_index == 4498 || pixel_index == 4500 || pixel_index == 4506 || ((pixel_index >= 4508) && (pixel_index <= 4510)) || pixel_index == 4512 || pixel_index == 4530 || pixel_index == 4584 || pixel_index == 4586 || pixel_index == 4588 || pixel_index == 4590 || ((pixel_index >= 4592) && (pixel_index <= 4593)) || ((pixel_index >= 4596) && (pixel_index <= 4601)) || ((pixel_index >= 4607) && (pixel_index <= 4608)) || ((pixel_index >= 4610) && (pixel_index <= 4611)) || ((pixel_index >= 4613) && (pixel_index <= 4614)) || pixel_index == 4616 || pixel_index == 4618 || ((pixel_index >= 4620) && (pixel_index <= 4621)) || ((pixel_index >= 4623) && (pixel_index <= 4625)) || ((pixel_index >= 4681) && (pixel_index <= 4682)) || pixel_index == 4684 || pixel_index == 4686 || pixel_index == 4688 || pixel_index == 4690 || pixel_index == 4692 || pixel_index == 4694 || ((pixel_index >= 4698) && (pixel_index <= 4704)) || pixel_index == 4706 || pixel_index == 4708 || pixel_index == 4712 || pixel_index == 4714 || pixel_index == 4716 || pixel_index == 4718 || pixel_index == 4782 || pixel_index == 4784 || pixel_index == 4786 || ((pixel_index >= 4788) && (pixel_index <= 4792)) || pixel_index == 4800 || pixel_index == 4802 || ((pixel_index >= 4804) && (pixel_index <= 4805)) || ((pixel_index >= 4807) && (pixel_index <= 4808)) || ((pixel_index >= 4810) && (pixel_index <= 4811)) || ((pixel_index >= 4813) && (pixel_index <= 4815)) || pixel_index == 4879 || pixel_index == 4881 || pixel_index == 4883 || ((pixel_index >= 4889) && (pixel_index <= 4896)) || pixel_index == 4902 || pixel_index == 4908 || pixel_index == 4910 || ((pixel_index >= 4976) && (pixel_index <= 4977)) || ((pixel_index >= 4979) && (pixel_index <= 4984)) || ((pixel_index >= 4992) && (pixel_index <= 4997)) || ((pixel_index >= 5000) && (pixel_index <= 5002)) || ((pixel_index >= 5004) && (pixel_index <= 5005)) || pixel_index == 5007 || pixel_index == 5072 || pixel_index == 5074 || pixel_index == 5078 || ((pixel_index >= 5080) && (pixel_index <= 5088)) || pixel_index == 5094 || pixel_index == 5102 || pixel_index == 5168 || ((pixel_index >= 5170) && (pixel_index <= 5175)) || pixel_index == 5179 || pixel_index == 5181 || ((pixel_index >= 5184) && (pixel_index <= 5189)) || pixel_index == 5192 || ((pixel_index >= 5194) && (pixel_index <= 5197)) || pixel_index == 5199 || ((pixel_index >= 5261) && (pixel_index <= 5262)) || ((pixel_index >= 5272) && (pixel_index <= 5278)) || pixel_index == 5280 || pixel_index == 5282 || pixel_index == 5284 || pixel_index == 5286 || pixel_index == 5290 || pixel_index == 5292 || pixel_index == 5294 || ((pixel_index >= 5354) && (pixel_index <= 5356)) || pixel_index == 5360 || ((pixel_index >= 5362) && (pixel_index <= 5365)) || ((pixel_index >= 5375) && (pixel_index <= 5377)) || ((pixel_index >= 5379) && (pixel_index <= 5380)) || pixel_index == 5382 || ((pixel_index >= 5384) && (pixel_index <= 5387)) || pixel_index == 5390 || ((pixel_index >= 5392) && (pixel_index <= 5393)) || ((pixel_index >= 5447) && (pixel_index <= 5450)) || pixel_index == 5452 || pixel_index == 5454 || ((pixel_index >= 5461) && (pixel_index <= 5462)) || ((pixel_index >= 5464) && (pixel_index <= 5469)) || pixel_index == 5472 || pixel_index == 5474 || pixel_index == 5478 || pixel_index == 5484 || pixel_index == 5486 || pixel_index == 5488 || pixel_index == 5490 || ((pixel_index >= 5541) && (pixel_index <= 5543)) || pixel_index == 5546 || pixel_index == 5551 || ((pixel_index >= 5553) && (pixel_index <= 5554)) || ((pixel_index >= 5567) && (pixel_index <= 5572)) || ((pixel_index >= 5574) && (pixel_index <= 5581)) || pixel_index == 5583 || pixel_index == 5585 || ((pixel_index >= 5588) && (pixel_index <= 5589)) || ((pixel_index >= 5592) && (pixel_index <= 5593)) || ((pixel_index >= 5595) && (pixel_index <= 5596)) || ((pixel_index >= 5598) && (pixel_index <= 5601)) || ((pixel_index >= 5603) && (pixel_index <= 5604)) || ((pixel_index >= 5606) && (pixel_index <= 5607)) || ((pixel_index >= 5609) && (pixel_index <= 5611)) || pixel_index == 5613 || pixel_index == 5615 || pixel_index == 5618 || ((pixel_index >= 5620) && (pixel_index <= 5624)) || ((pixel_index >= 5626) && (pixel_index <= 5627)) || ((pixel_index >= 5629) && (pixel_index <= 5637)) || pixel_index == 5639 || pixel_index == 5642 || pixel_index == 5644 || pixel_index == 5646 || pixel_index == 5648 || pixel_index == 5650 || pixel_index == 5652 || pixel_index == 5654 || ((pixel_index >= 5656) && (pixel_index <= 5662)) || pixel_index == 5664 || pixel_index == 5666 || pixel_index == 5668 || ((pixel_index >= 5682) && (pixel_index <= 5683)) || pixel_index == 5687 || pixel_index == 5689 || ((pixel_index >= 5692) && (pixel_index <= 5694)) || pixel_index == 5696 || pixel_index == 5698 || pixel_index == 5700 || pixel_index == 5703 || pixel_index == 5705 || pixel_index == 5707 || pixel_index == 5709 || pixel_index == 5718 || pixel_index == 5720 || pixel_index == 5722 || ((pixel_index >= 5733) && (pixel_index <= 5735)) || pixel_index == 5737 || pixel_index == 5739 || ((pixel_index >= 5741) && (pixel_index <= 5742)) || pixel_index == 5744 || pixel_index == 5749 || pixel_index == 5751 || ((pixel_index >= 5759) && (pixel_index <= 5763)) || ((pixel_index >= 5766) && (pixel_index <= 5774)) || pixel_index == 5776 || ((pixel_index >= 5780) && (pixel_index <= 5783)) || pixel_index == 5785 || pixel_index == 5791 || pixel_index == 5793 || pixel_index == 5796 || ((pixel_index >= 5802) && (pixel_index <= 5803)) || ((pixel_index >= 5806) && (pixel_index <= 5807)) || ((pixel_index >= 5809) && (pixel_index <= 5812)) || ((pixel_index >= 5814) && (pixel_index <= 5815)) || ((pixel_index >= 5817) && (pixel_index <= 5825)) || pixel_index == 5827 || ((pixel_index >= 5834) && (pixel_index <= 5835)) || pixel_index == 5838 || pixel_index == 5840 || ((pixel_index >= 5842) && (pixel_index <= 5845)) || ((pixel_index >= 5847) && (pixel_index <= 5850)) || ((pixel_index >= 5852) && (pixel_index <= 5853)) || pixel_index == 5856 || pixel_index == 5860 || pixel_index == 5872 || pixel_index == 5875 || pixel_index == 5882 || ((pixel_index >= 5884) && (pixel_index <= 5885)) || pixel_index == 5891 || pixel_index == 5893 || pixel_index == 5895 || pixel_index == 5897 || pixel_index == 5900 || pixel_index == 5905 || pixel_index == 5907 || pixel_index == 5909 || pixel_index == 5911 || ((pixel_index >= 5925) && (pixel_index <= 5929)) || ((pixel_index >= 5932) && (pixel_index <= 5933)) || pixel_index == 5935 || pixel_index == 5939 || pixel_index == 5941 || pixel_index == 5943 || pixel_index == 5945 || pixel_index == 5949 || ((pixel_index >= 5952) && (pixel_index <= 5953)) || pixel_index == 5955 || ((pixel_index >= 5957) && (pixel_index <= 5964)) || ((pixel_index >= 5966) && (pixel_index <= 5967)) || pixel_index == 5969 || ((pixel_index >= 5972) && (pixel_index <= 5974)) || ((pixel_index >= 5976) && (pixel_index <= 5977)) || ((pixel_index >= 5982) && (pixel_index <= 5983)) || pixel_index == 5985 || pixel_index == 5988 || pixel_index == 5991 || ((pixel_index >= 5993) && (pixel_index <= 5994)) || ((pixel_index >= 5997) && (pixel_index <= 5999)) || ((pixel_index >= 6001) && (pixel_index <= 6002)) || pixel_index == 6004 || ((pixel_index >= 6007) && (pixel_index <= 6016)) || ((pixel_index >= 6018) && (pixel_index <= 6019)) || pixel_index == 6021 || ((pixel_index >= 6025) && (pixel_index <= 6026)) || pixel_index == 6031 || ((pixel_index >= 6033) && (pixel_index <= 6037)) || ((pixel_index >= 6039) && (pixel_index <= 6043)) || ((pixel_index >= 6045) && (pixel_index <= 6048)) || pixel_index == 6050 || pixel_index == 6052 || pixel_index == 6064 || pixel_index == 6066 || pixel_index == 6068 || pixel_index == 6070 || ((pixel_index >= 6074) && (pixel_index <= 6075)) || pixel_index == 6081 || pixel_index == 6083 || pixel_index == 6085 || pixel_index == 6087 || pixel_index == 6089 || ((pixel_index >= 6091) && (pixel_index <= 6092)) || pixel_index == 6116 || ((pixel_index >= 6118) && (pixel_index <= 6120)) || ((pixel_index >= 6122) && (pixel_index <= 6125)) || pixel_index == 6127) oled_data = 16'b0101001101010001;
    else if (pixel_index == 97 || pixel_index == 99 || pixel_index == 101 || pixel_index == 103 || pixel_index == 105 || pixel_index == 107 || pixel_index == 109 || pixel_index == 111 || pixel_index == 113 || pixel_index == 115 || pixel_index == 117 || pixel_index == 119 || pixel_index == 121 || pixel_index == 123 || pixel_index == 125 || pixel_index == 127 || pixel_index == 129 || pixel_index == 131 || pixel_index == 133 || pixel_index == 135 || pixel_index == 137 || pixel_index == 139 || pixel_index == 141 || pixel_index == 143 || pixel_index == 145 || pixel_index == 147 || pixel_index == 149 || pixel_index == 151 || pixel_index == 153 || pixel_index == 155 || pixel_index == 157 || pixel_index == 159 || pixel_index == 161 || pixel_index == 163 || pixel_index == 165 || pixel_index == 167 || pixel_index == 169 || pixel_index == 171 || pixel_index == 173 || pixel_index == 175 || pixel_index == 177 || pixel_index == 179 || pixel_index == 181 || pixel_index == 183 || pixel_index == 185 || pixel_index == 187 || pixel_index == 189 || pixel_index == 347 || pixel_index == 481 || pixel_index == 483 || pixel_index == 485 || pixel_index == 487 || pixel_index == 497 || pixel_index == 499 || pixel_index == 509 || pixel_index == 511 || pixel_index == 523 || pixel_index == 673 || pixel_index == 733 || pixel_index == 865 || pixel_index == 867 || pixel_index == 875 || pixel_index == 877 || pixel_index == 881 || pixel_index == 1079 || pixel_index == 1123 || pixel_index == 1249 || pixel_index == 1251 || pixel_index == 1313 || pixel_index == 1331 || pixel_index == 1441 || pixel_index == 1453 || pixel_index == 1459 || pixel_index == 1633 || pixel_index == 1649 || pixel_index == 1651 || pixel_index == 1655 || pixel_index == 1707 || pixel_index == 1709 || pixel_index == 1713 || pixel_index == 1756 || pixel_index == 1833 || pixel_index == 1911 || pixel_index == 2017 || pixel_index == 2033 || pixel_index == 2035 || pixel_index == 2294 || pixel_index == 2474 || pixel_index == 2476 || pixel_index == 2597 || pixel_index == 2599 || pixel_index == 2609 || pixel_index == 2667 || pixel_index == 2787 || pixel_index == 2789 || pixel_index == 2799 || pixel_index == 2801 || pixel_index == 3046 || pixel_index == 3171 || pixel_index == 3237 || pixel_index == 3369 || pixel_index == 3381 || pixel_index == 3561 || pixel_index == 3751 || pixel_index == 3753 || pixel_index == 4311 || pixel_index == 4337 || pixel_index == 4483 || pixel_index == 4693 || pixel_index == 4719 || pixel_index == 5079 || pixel_index == 5180 || pixel_index == 5281 || pixel_index == 5283 || pixel_index == 5291 || pixel_index == 5473 || pixel_index == 5665 || pixel_index == 5667 || pixel_index == 5719 || pixel_index == 5906 || pixel_index == 5940 || pixel_index == 5944 || pixel_index == 6049 || pixel_index == 6069 || pixel_index == 6090 || pixel_index == 6121) oled_data = 16'b0101101110010010;
    else if (pixel_index == 191 || pixel_index == 289 || pixel_index == 291 || pixel_index == 345 || pixel_index == 540 || pixel_index == 542 || pixel_index == 546 || pixel_index == 548 || pixel_index == 550 || pixel_index == 558 || pixel_index == 560 || pixel_index == 562 || pixel_index == 570 || pixel_index == 572 || pixel_index == 675 || pixel_index == 677 || pixel_index == 731 || pixel_index == 814 || pixel_index == 1057 || pixel_index == 1059 || pixel_index == 1071 || pixel_index == 1077 || pixel_index == 1081 || pixel_index == 1119 || pixel_index == 1121 || pixel_index == 1257 || pixel_index == 1259 || pixel_index == 1261 || pixel_index == 1263 || pixel_index == 1267 || pixel_index == 1269 || pixel_index == 1271 || pixel_index == 1311 || pixel_index == 1443 || pixel_index == 1449 || pixel_index == 1451 || pixel_index == 1455 || pixel_index == 1461 || pixel_index == 1463 || pixel_index == 1502 || pixel_index == 1504 || pixel_index == 1530 || pixel_index == 1582 || pixel_index == 1639 || pixel_index == 1641 || pixel_index == 1643 || pixel_index == 1645 || pixel_index == 1653 || pixel_index == 1699 || pixel_index == 1701 || pixel_index == 1711 || pixel_index == 1825 || pixel_index == 1829 || pixel_index == 1831 || pixel_index == 1835 || pixel_index == 1837 || pixel_index == 1887 || pixel_index == 1919 || pixel_index == 1946 || pixel_index == 1948 || pixel_index == 2021 || pixel_index == 2023 || pixel_index == 2025 || pixel_index == 2078 || pixel_index == 2102 || pixel_index == 2110 || pixel_index == 2211 || pixel_index == 2213 || pixel_index == 2215 || pixel_index == 2217 || pixel_index == 2219 || pixel_index == 2595 || pixel_index == 2607 || pixel_index == 2665 || pixel_index == 2797 || pixel_index == 3164 || pixel_index == 3181 || pixel_index == 3183 || pixel_index == 3191 || pixel_index == 3383 || pixel_index == 3432 || pixel_index == 3434 || pixel_index == 3547 || pixel_index == 3740 || pixel_index == 3742 || pixel_index == 3755 || pixel_index == 3757 || pixel_index == 3955 || pixel_index == 3957 || pixel_index == 4016 || pixel_index == 4018 || pixel_index == 4119 || pixel_index == 4147 || pixel_index == 4149 || pixel_index == 4202 || pixel_index == 4290 || pixel_index == 4339 || pixel_index == 4343 || pixel_index == 4501 || pixel_index == 4503 || pixel_index == 4505 || pixel_index == 4529 || pixel_index == 4585 || pixel_index == 4587 || pixel_index == 4589 || pixel_index == 4604 || pixel_index == 4606 || pixel_index == 4691 || pixel_index == 4695 || pixel_index == 4697 || pixel_index == 4707 || pixel_index == 4709 || pixel_index == 4713 || pixel_index == 4715 || pixel_index == 4882 || pixel_index == 4884 || pixel_index == 4886 || pixel_index == 4888 || pixel_index == 4909 || pixel_index == 4911 || pixel_index == 5073 || pixel_index == 5075 || pixel_index == 5077 || pixel_index == 5089 || pixel_index == 5091 || pixel_index == 5093 || pixel_index == 5101 || pixel_index == 5176 || pixel_index == 5178 || pixel_index == 5182 || pixel_index == 5285 || pixel_index == 5289 || pixel_index == 5295 || pixel_index == 5451 || pixel_index == 5485 || pixel_index == 5487 || pixel_index == 5489 || pixel_index == 5597 || pixel_index == 5638 || pixel_index == 5647 || pixel_index == 5649 || pixel_index == 5695 || pixel_index == 5697 || pixel_index == 5706 || pixel_index == 5717 || pixel_index == 5723 || pixel_index == 5740 || pixel_index == 5748 || pixel_index == 5750 || pixel_index == 5752 || pixel_index == 5754 || pixel_index == 5756 || pixel_index == 5789 || pixel_index == 5833 || pixel_index == 5837 || pixel_index == 5839 || pixel_index == 5857 || pixel_index == 5881 || pixel_index == 5892 || pixel_index == 5898 || pixel_index == 5902 || pixel_index == 5908 || pixel_index == 5910 || pixel_index == 5938 || pixel_index == 5942 || pixel_index == 5946 || pixel_index == 6020 || pixel_index == 6022 || pixel_index == 6024 || pixel_index == 6065 || pixel_index == 6073 || pixel_index == 6084) oled_data = 16'b0101001110010010;
    else if (pixel_index == 196 || pixel_index == 202 || pixel_index == 208 || pixel_index == 214 || pixel_index == 220 || pixel_index == 226 || pixel_index == 232 || pixel_index == 238 || pixel_index == 252 || pixel_index == 258 || pixel_index == 264 || pixel_index == 270 || pixel_index == 276 || pixel_index == 282 || pixel_index == 294 || pixel_index == 300 || pixel_index == 306 || pixel_index == 312 || pixel_index == 318 || pixel_index == 332 || pixel_index == 352 || pixel_index == 358 || pixel_index == 364 || pixel_index == 370 || pixel_index == 376 || pixel_index == 382 || pixel_index == 393 || pixel_index == 399 || pixel_index == 405 || pixel_index == 411 || pixel_index == 429 || pixel_index == 449 || pixel_index == 455 || pixel_index == 461 || pixel_index == 467 || pixel_index == 473 || pixel_index == 479 || pixel_index == 490 || pixel_index == 492 || pixel_index == 494 || pixel_index == 502 || pixel_index == 504 || pixel_index == 506 || pixel_index == 584 || pixel_index == 592 || pixel_index == 596 || pixel_index == 604 || pixel_index == 621 || pixel_index == 639 || pixel_index == 648 || pixel_index == 652 || pixel_index == 660 || pixel_index == 664 || pixel_index == 671 || pixel_index == 684 || pixel_index == 686 || pixel_index == 690 || pixel_index == 696 || pixel_index == 698 || pixel_index == 702 || pixel_index == 738 || pixel_index == 740 || pixel_index == 746 || pixel_index == 750 || pixel_index == 752 || pixel_index == 758 || pixel_index == 762 || pixel_index == 772 || pixel_index == 775 || pixel_index == 777 || pixel_index == 784 || pixel_index == 788 || pixel_index == 796 || pixel_index == 812 || pixel_index == 830 || pixel_index == 839 || pixel_index == 844 || pixel_index == 852 || pixel_index == 856 || pixel_index == 859 || pixel_index == 863 || pixel_index == 886 || pixel_index == 888 || pixel_index == 890 || pixel_index == 928 || pixel_index == 930 || pixel_index == 932 || pixel_index == 936 || pixel_index == 938 || pixel_index == 942 || pixel_index == 944 || pixel_index == 946 || pixel_index == 950 || pixel_index == 965 || pixel_index == 967 || pixel_index == 969 || pixel_index == 974 || pixel_index == 978 || pixel_index == 980 || pixel_index == 987 || pixel_index == 1005 || pixel_index == 1020 || pixel_index == 1022 || pixel_index == 1029 || pixel_index == 1035 || pixel_index == 1043 || pixel_index == 1047 || pixel_index == 1049 || pixel_index == 1051 || pixel_index == 1053 || pixel_index == 1055 || pixel_index == 1066 || pixel_index == 1068 || pixel_index == 1128 || pixel_index == 1134 || pixel_index == 1136 || pixel_index == 1140 || pixel_index == 1156 || pixel_index == 1158 || pixel_index == 1160 || pixel_index == 1168 || pixel_index == 1170 || pixel_index == 1178 || pixel_index == 1196 || pixel_index == 1213 || pixel_index == 1220 || pixel_index == 1225 || pixel_index == 1233 || pixel_index == 1237 || pixel_index == 1239 || pixel_index == 1241 || pixel_index == 1243 || pixel_index == 1247 || pixel_index == 1318 || pixel_index == 1322 || pixel_index == 1324 || pixel_index == 1326 || pixel_index == 1328 || pixel_index == 1349 || pixel_index == 1351 || pixel_index == 1361 || pixel_index == 1368 || pixel_index == 1370 || pixel_index == 1390 || pixel_index == 1405 || pixel_index == 1410 || pixel_index == 1412 || pixel_index == 1415 || pixel_index == 1417 || pixel_index == 1426 || pixel_index == 1429 || pixel_index == 1431 || pixel_index == 1433 || pixel_index == 1435 || pixel_index == 1439 || pixel_index == 1469 || pixel_index == 1509 || pixel_index == 1515 || pixel_index == 1519 || pixel_index == 1521 || pixel_index == 1540 || pixel_index == 1542 || pixel_index == 1552 || pixel_index == 1561 || pixel_index == 1596 || pixel_index == 1602 || pixel_index == 1607 || pixel_index == 1619 || pixel_index == 1623 || pixel_index == 1625 || pixel_index == 1628 || pixel_index == 1630 || pixel_index == 1661 || pixel_index == 1694 || pixel_index == 1730 || pixel_index == 1732 || pixel_index == 1752 || pixel_index == 1754 || pixel_index == 1789 || pixel_index == 1794 || pixel_index == 1798 || pixel_index == 1802 || pixel_index == 1810 || pixel_index == 1812 || pixel_index == 1814 || pixel_index == 1816 || pixel_index == 1818 || pixel_index == 1820 || pixel_index == 1822 || pixel_index == 1842 || pixel_index == 1844 || pixel_index == 1846 || pixel_index == 1892 || pixel_index == 1900 || pixel_index == 1902 || pixel_index == 1904 || pixel_index == 1923 || pixel_index == 1930 || pixel_index == 1935 || pixel_index == 1941 || pixel_index == 1944 || pixel_index == 1951 || pixel_index == 1980 || pixel_index == 1986 || pixel_index == 1990 || pixel_index == 1994 || pixel_index == 2003 || pixel_index == 2005 || pixel_index == 2013 || pixel_index == 2028 || pixel_index == 2083 || pixel_index == 2095 || pixel_index == 2114 || pixel_index == 2125 || pixel_index == 2127 || pixel_index == 2132 || pixel_index == 2134 || pixel_index == 2136 || pixel_index == 2138 || pixel_index == 2173 || pixel_index == 2180 || pixel_index == 2182 || pixel_index == 2184 || pixel_index == 2192 || pixel_index == 2194 || pixel_index == 2196 || pixel_index == 2200 || pixel_index == 2202 || pixel_index == 2204 || pixel_index == 2224 || pixel_index == 2273 || pixel_index == 2281 || pixel_index == 2285 || pixel_index == 2301 || pixel_index == 2303 || pixel_index == 2305 || pixel_index == 2316 || pixel_index == 2318 || pixel_index == 2328 || pixel_index == 2330 || pixel_index == 2367 || pixel_index == 2370 || pixel_index == 2372 || pixel_index == 2374 || pixel_index == 2382 || pixel_index == 2384 || pixel_index == 2386 || pixel_index == 2388 || pixel_index == 2391 || pixel_index == 2393 || pixel_index == 2395 || pixel_index == 2402 || pixel_index == 2404 || pixel_index == 2406 || pixel_index == 2410 || pixel_index == 2416 || pixel_index == 2418 || pixel_index == 2485 || pixel_index == 2492 || pixel_index == 2497 || pixel_index == 2505 || pixel_index == 2508 || pixel_index == 2510 || pixel_index == 2517 || pixel_index == 2519 || pixel_index == 2521 || pixel_index == 2562 || pixel_index == 2564 || pixel_index == 2566 || pixel_index == 2573 || pixel_index == 2575 || pixel_index == 2577 || pixel_index == 2579 || pixel_index == 2583 || pixel_index == 2682 || pixel_index == 2684 || pixel_index == 2686 || pixel_index == 2689 || pixel_index == 2696 || pixel_index == 2698 || pixel_index == 2709 || pixel_index == 2711 || pixel_index == 2754 || pixel_index == 2756 || pixel_index == 2758 || pixel_index == 2760 || pixel_index == 2765 || pixel_index == 2767 || pixel_index == 2769 || pixel_index == 2773 || pixel_index == 2775 || pixel_index == 2858 || pixel_index == 2866 || pixel_index == 2872 || pixel_index == 2876 || pixel_index == 2878 || pixel_index == 2881 || pixel_index == 2886 || pixel_index == 2888 || pixel_index == 2890 || pixel_index == 2892 || pixel_index == 2898 || pixel_index == 2902 || pixel_index == 2947 || pixel_index == 2949 || pixel_index == 2951 || pixel_index == 2955 || pixel_index == 2957 || pixel_index == 2964 || pixel_index == 2966 || pixel_index == 2978 || pixel_index == 2990 || pixel_index == 2992 || pixel_index == 3049 || pixel_index == 3059 || pixel_index == 3063 || pixel_index == 3065 || pixel_index == 3073 || pixel_index == 3078 || pixel_index == 3080 || pixel_index == 3082 || pixel_index == 3090 || pixel_index == 3094 || pixel_index == 3138 || pixel_index == 3140 || pixel_index == 3147 || pixel_index == 3149 || pixel_index == 3151 || pixel_index == 3153 || pixel_index == 3157 || pixel_index == 3250 || pixel_index == 3256 || pixel_index == 3258 || pixel_index == 3262 || pixel_index == 3265 || pixel_index == 3268 || pixel_index == 3270 || pixel_index == 3272 || pixel_index == 3274 || pixel_index == 3276 || pixel_index == 3280 || pixel_index == 3282 || pixel_index == 3284 || pixel_index == 3331 || pixel_index == 3340 || pixel_index == 3342 || pixel_index == 3347 || pixel_index == 3355 || pixel_index == 3359 || pixel_index == 3374 || pixel_index == 3441 || pixel_index == 3445 || pixel_index == 3447 || pixel_index == 3449 || pixel_index == 3457 || pixel_index == 3459 || pixel_index == 3461 || pixel_index == 3463 || pixel_index == 3472 || pixel_index == 3474 || pixel_index == 3476 || pixel_index == 3523 || pixel_index == 3526 || pixel_index == 3531 || pixel_index == 3533 || pixel_index == 3535 || pixel_index == 3550 || pixel_index == 3564 || pixel_index == 3574 || pixel_index == 3620 || pixel_index == 3624 || pixel_index == 3632 || pixel_index == 3636 || pixel_index == 3638 || pixel_index == 3640 || pixel_index == 3649 || pixel_index == 3653 || pixel_index == 3663 || pixel_index == 3665 || pixel_index == 3667 || pixel_index == 3714 || pixel_index == 3718 || pixel_index == 3721 || pixel_index == 3723 || pixel_index == 3725 || pixel_index == 3766 || pixel_index == 3812 || pixel_index == 3822 || pixel_index == 3826 || pixel_index == 3828 || pixel_index == 3830 || pixel_index == 3832 || pixel_index == 3834 || pixel_index == 3839 || pixel_index == 3841 || pixel_index == 3845 || pixel_index == 3854 || pixel_index == 3856 || pixel_index == 3858 || pixel_index == 3907 || pixel_index == 3910 || pixel_index == 3912 || pixel_index == 3914 || pixel_index == 3919 || pixel_index == 3931 || pixel_index == 3933 || pixel_index == 3938 || pixel_index == 3944 || pixel_index == 3946 || pixel_index == 3948 || pixel_index == 4013 || pixel_index == 4024 || pixel_index == 4031 || pixel_index == 4033 || pixel_index == 4045 || pixel_index == 4047 || pixel_index == 4049 || pixel_index == 4055 || pixel_index == 4099 || pixel_index == 4101 || pixel_index == 4103 || pixel_index == 4105 || pixel_index == 4107 || pixel_index == 4124 || pixel_index == 4138 || pixel_index == 4140 || pixel_index == 4153 || pixel_index == 4205 || pixel_index == 4207 || pixel_index == 4209 || pixel_index == 4211 || pixel_index == 4217 || pixel_index == 4221 || pixel_index == 4223 || pixel_index == 4225 || pixel_index == 4227 || pixel_index == 4238 || pixel_index == 4240 || pixel_index == 4292 || pixel_index == 4294 || pixel_index == 4296 || pixel_index == 4308 || pixel_index == 4314 || pixel_index == 4324 || pixel_index == 4326 || pixel_index == 4328 || pixel_index == 4330 || pixel_index == 4332 || pixel_index == 4393 || pixel_index == 4395 || pixel_index == 4397 || pixel_index == 4399 || pixel_index == 4401 || pixel_index == 4403 || pixel_index == 4411 || pixel_index == 4415 || pixel_index == 4417 || pixel_index == 4429 || pixel_index == 4431 || pixel_index == 4436 || pixel_index == 4485 || pixel_index == 4487 || pixel_index == 4496 || pixel_index == 4514 || pixel_index == 4516 || pixel_index == 4518 || pixel_index == 4520 || pixel_index == 4522 || pixel_index == 4524 || pixel_index == 4591 || pixel_index == 4594 || pixel_index == 4602 || pixel_index == 4609 || pixel_index == 4622 || pixel_index == 4779 || pixel_index == 4781 || pixel_index == 4783 || pixel_index == 4785 || pixel_index == 4797 || pixel_index == 4799 || pixel_index == 4801 || pixel_index == 4806 || pixel_index == 4898 || pixel_index == 4900 || pixel_index == 4906 || pixel_index == 4975 || pixel_index == 4985 || pixel_index == 4987 || pixel_index == 4989 || pixel_index == 4991 || pixel_index == 4998 || pixel_index == 5096 || pixel_index == 5098 || pixel_index == 5191 || pixel_index == 5264 || pixel_index == 5266 || pixel_index == 5268 || pixel_index == 5270 || pixel_index == 5279 || pixel_index == 5358 || pixel_index == 5367 || pixel_index == 5378 || pixel_index == 5383 || pixel_index == 5388 || pixel_index == 5456 || pixel_index == 5458 || pixel_index == 5470 || pixel_index == 5480 || pixel_index == 5482 || pixel_index == 5544 || pixel_index == 5548 || pixel_index == 5550 || pixel_index == 5557 || pixel_index == 5559 || pixel_index == 5561 || pixel_index == 5563 || pixel_index == 5573 || pixel_index == 5591 || pixel_index == 5594 || pixel_index == 5602 || pixel_index == 5605 || pixel_index == 5614 || pixel_index == 5617 || pixel_index == 5625 || pixel_index == 5628 || pixel_index == 5641 || pixel_index == 5651 || pixel_index == 5663 || pixel_index == 5672 || pixel_index == 5674 || pixel_index == 5678 || pixel_index == 5680 || pixel_index == 5684 || pixel_index == 5686 || pixel_index == 5691 || pixel_index == 5702 || pixel_index == 5704 || pixel_index == 5712 || pixel_index == 5715 || pixel_index == 5730 || pixel_index == 5764 || pixel_index == 5777 || pixel_index == 5784 || pixel_index == 5795 || pixel_index == 5805 || pixel_index == 5816 || pixel_index == 5829 || pixel_index == 5831 || pixel_index == 5841 || pixel_index == 5851 || pixel_index == 5854 || pixel_index == 5862 || pixel_index == 5864 || pixel_index == 5866 || pixel_index == 5868 || pixel_index == 5870 || pixel_index == 5874 || pixel_index == 5883 || pixel_index == 5887 || pixel_index == 5889 || pixel_index == 5894 || pixel_index == 5896 || pixel_index == 5904 || pixel_index == 5913 || pixel_index == 5915 || pixel_index == 5917 || pixel_index == 5921 || pixel_index == 5923 || pixel_index == 5931 || pixel_index == 5951 || pixel_index == 5954 || pixel_index == 5965 || pixel_index == 5975 || pixel_index == 5980 || pixel_index == 5986 || pixel_index == 5995 || pixel_index == 6005 || pixel_index == 6030 || pixel_index == 6032 || pixel_index == 6044 || pixel_index == 6056 || pixel_index == 6058 || pixel_index == 6067 || pixel_index == 6077 || pixel_index == 6079 || pixel_index == 6086 || pixel_index == 6088 || pixel_index == 6095 || pixel_index == 6097 || pixel_index == 6099 || pixel_index == 6103 || pixel_index == 6107 || pixel_index == 6109 || pixel_index == 6111 || pixel_index == 6113 || pixel_index == 6129 || pixel_index == 6131 || pixel_index == 6133 || pixel_index == 6135 || pixel_index == 6143) oled_data = 16'b0101001101010010;
    else if (pixel_index == 287 || pixel_index == 290 || pixel_index == 478 || pixel_index == 539 || pixel_index == 541 || pixel_index == 543 || pixel_index == 545 || pixel_index == 547 || pixel_index == 549 || pixel_index == 551 || pixel_index == 557 || pixel_index == 559 || pixel_index == 561 || pixel_index == 563 || pixel_index == 569 || pixel_index == 571 || pixel_index == 676 || pixel_index == 688 || pixel_index == 700 || pixel_index == 717 || pixel_index == 748 || pixel_index == 760 || pixel_index == 1054 || pixel_index == 1058 || pixel_index == 1064 || pixel_index == 1070 || pixel_index == 1076 || pixel_index == 1082 || pixel_index == 1120 || pixel_index == 1138 || pixel_index == 1144 || pixel_index == 1159 || pixel_index == 1215 || pixel_index == 1258 || pixel_index == 1260 || pixel_index == 1262 || pixel_index == 1264 || pixel_index == 1266 || pixel_index == 1268 || pixel_index == 1270 || pixel_index == 1272 || pixel_index == 1274 || pixel_index == 1352 || pixel_index == 1444 || pixel_index == 1446 || pixel_index == 1450 || pixel_index == 1456 || pixel_index == 1462 || pixel_index == 1501 || pixel_index == 1503 || pixel_index == 1505 || pixel_index == 1511 || pixel_index == 1523 || pixel_index == 1529 || pixel_index == 1551 || pixel_index == 1557 || pixel_index == 1615 || pixel_index == 1627 || pixel_index == 1629 || pixel_index == 1638 || pixel_index == 1640 || pixel_index == 1642 || pixel_index == 1644 || pixel_index == 1678 || pixel_index == 1698 || pixel_index == 1700 || pixel_index == 1702 || pixel_index == 1791 || pixel_index == 1819 || pixel_index == 1826 || pixel_index == 1828 || pixel_index == 1830 || pixel_index == 1836 || pixel_index == 1848 || pixel_index == 1850 || pixel_index == 1894 || pixel_index == 1898 || pixel_index == 1906 || pixel_index == 1931 || pixel_index == 1943 || pixel_index == 2015 || pixel_index == 2022 || pixel_index == 2024 || pixel_index == 2043 || pixel_index == 2047 || pixel_index == 2077 || pixel_index == 2099 || pixel_index == 2101 || pixel_index == 2109 || pixel_index == 2122 || pixel_index == 2133 || pixel_index == 2135 || pixel_index == 2137 || pixel_index == 2174 || pixel_index == 2185 || pixel_index == 2191 || pixel_index == 2193 || pixel_index == 2203 || pixel_index == 2212 || pixel_index == 2214 || pixel_index == 2216 || pixel_index == 2220 || pixel_index == 2275 || pixel_index == 2297 || pixel_index == 2314 || pixel_index == 2329 || pixel_index == 2368 || pixel_index == 2385 || pixel_index == 2392 || pixel_index == 2396 || pixel_index == 2483 || pixel_index == 2486 || pixel_index == 2507 || pixel_index == 2518 || pixel_index == 2520 || pixel_index == 2576 || pixel_index == 2587 || pixel_index == 2594 || pixel_index == 2606 || pixel_index == 2662 || pixel_index == 2670 || pixel_index == 2674 || pixel_index == 2678 || pixel_index == 2685 || pixel_index == 2761 || pixel_index == 2768 || pixel_index == 2776 || pixel_index == 2779 || pixel_index == 2783 || pixel_index == 2792 || pixel_index == 2806 || pixel_index == 2850 || pixel_index == 2852 || pixel_index == 2854 || pixel_index == 2870 || pixel_index == 2893 || pixel_index == 2952 || pixel_index == 2968 || pixel_index == 2982 || pixel_index == 2984 || pixel_index == 2986 || pixel_index == 2994 || pixel_index == 3043 || pixel_index == 3053 || pixel_index == 3152 || pixel_index == 3155 || pixel_index == 3161 || pixel_index == 3165 || pixel_index == 3174 || pixel_index == 3182 || pixel_index == 3184 || pixel_index == 3186 || pixel_index == 3190 || pixel_index == 3244 || pixel_index == 3246 || pixel_index == 3259 || pixel_index == 3269 || pixel_index == 3275 || pixel_index == 3346 || pixel_index == 3349 || pixel_index == 3362 || pixel_index == 3376 || pixel_index == 3433 || pixel_index == 3450 || pixel_index == 3460 || pixel_index == 3479 || pixel_index == 3527 || pixel_index == 3534 || pixel_index == 3536 || pixel_index == 3541 || pixel_index == 3544 || pixel_index == 3568 || pixel_index == 3570 || pixel_index == 3572 || pixel_index == 3626 || pixel_index == 3628 || pixel_index == 3644 || pixel_index == 3647 || pixel_index == 3660 || pixel_index == 3670 || pixel_index == 3720 || pixel_index == 3726 || pixel_index == 3731 || pixel_index == 3758 || pixel_index == 3814 || pixel_index == 3818 || pixel_index == 3829 || pixel_index == 3835 || pixel_index == 3837 || pixel_index == 3851 || pixel_index == 3859 || pixel_index == 3909 || pixel_index == 3918 || pixel_index == 3920 || pixel_index == 3922 || pixel_index == 3935 || pixel_index == 4003 || pixel_index == 4029 || pixel_index == 4043 || pixel_index == 4052 || pixel_index == 4054 || pixel_index == 4102 || pixel_index == 4108 || pixel_index == 4111 || pixel_index == 4114 || pixel_index == 4130 || pixel_index == 4142 || pixel_index == 4152 || pixel_index == 4216 || pixel_index == 4218 || pixel_index == 4220 || pixel_index == 4222 || pixel_index == 4228 || pixel_index == 4234 || pixel_index == 4236 || pixel_index == 4243 || pixel_index == 4291 || pixel_index == 4298 || pixel_index == 4300 || pixel_index == 4302 || pixel_index == 4304 || pixel_index == 4306 || pixel_index == 4389 || pixel_index == 4391 || pixel_index == 4404 || pixel_index == 4410 || pixel_index == 4419 || pixel_index == 4421 || pixel_index == 4425 || pixel_index == 4428 || pixel_index == 4435 || pixel_index == 4489 || pixel_index == 4491 || pixel_index == 4494 || pixel_index == 4502 || pixel_index == 4504 || pixel_index == 4511 || pixel_index == 4526 || pixel_index == 4528 || pixel_index == 4595 || pixel_index == 4603 || pixel_index == 4605 || pixel_index == 4612 || pixel_index == 4617 || pixel_index == 4619 || pixel_index == 4683 || pixel_index == 4685 || pixel_index == 4696 || pixel_index == 4710 || pixel_index == 4787 || pixel_index == 4793 || pixel_index == 4803 || pixel_index == 4809 || pixel_index == 4877 || pixel_index == 4885 || pixel_index == 4887 || pixel_index == 4978 || pixel_index == 4999 || pixel_index == 5006 || pixel_index == 5076 || pixel_index == 5090 || pixel_index == 5092 || pixel_index == 5100 || pixel_index == 5169 || pixel_index == 5177 || pixel_index == 5183 || pixel_index == 5190 || pixel_index == 5193 || pixel_index == 5271 || pixel_index == 5288 || pixel_index == 5359 || pixel_index == 5361 || pixel_index == 5381 || pixel_index == 5389 || pixel_index == 5391 || pixel_index == 5453 || pixel_index == 5463 || pixel_index == 5471 || pixel_index == 5547 || pixel_index == 5552 || pixel_index == 5555 || pixel_index == 5582 || pixel_index == 5584 || pixel_index == 5640 || pixel_index == 5645 || pixel_index == 5653 || pixel_index == 5655 || pixel_index == 5711 || pixel_index == 5713 || pixel_index == 5716 || pixel_index == 5724 || pixel_index == 5743 || pixel_index == 5745 || pixel_index == 5747 || pixel_index == 5753 || pixel_index == 5755 || pixel_index == 5757 || pixel_index == 5765 || pixel_index == 5775 || pixel_index == 5778 || pixel_index == 5786 || pixel_index == 5788 || pixel_index == 5790 || pixel_index == 5792 || pixel_index == 5794 || pixel_index == 5797 || pixel_index == 5799 || pixel_index == 5801 || pixel_index == 5813 || pixel_index == 5826 || pixel_index == 5832 || pixel_index == 5836 || pixel_index == 5846 || pixel_index == 5855 || pixel_index == 5858 || pixel_index == 5880 || pixel_index == 5899 || pixel_index == 5901 || pixel_index == 5903 || pixel_index == 5924 || pixel_index == 5934 || pixel_index == 5937 || pixel_index == 5947 || pixel_index == 5970 || pixel_index == 5978 || pixel_index == 5981 || pixel_index == 5984 || pixel_index == 5987 || pixel_index == 5989 || pixel_index == 6003 || pixel_index == 6006 || pixel_index == 6017 || pixel_index == 6023 || pixel_index == 6038 || pixel_index == 6062 || pixel_index == 6072 || pixel_index == 6096 || pixel_index == 6101 || pixel_index == 6117 || pixel_index == 6139) oled_data = 16'b0101101101010001;
    else if (pixel_index == 293 || pixel_index == 299 || pixel_index == 305 || pixel_index == 311 || pixel_index == 317 || pixel_index == 333 || pixel_index == 353 || pixel_index == 359 || pixel_index == 365 || pixel_index == 371 || pixel_index == 377 || pixel_index == 489 || pixel_index == 491 || pixel_index == 493 || pixel_index == 495 || pixel_index == 501 || pixel_index == 503 || pixel_index == 505 || pixel_index == 507 || pixel_index == 525 || pixel_index == 679 || pixel_index == 685 || pixel_index == 691 || pixel_index == 697 || pixel_index == 739 || pixel_index == 745 || pixel_index == 751 || pixel_index == 757 || pixel_index == 763 || pixel_index == 767 || pixel_index == 798 || pixel_index == 869 || pixel_index == 871 || pixel_index == 873 || pixel_index == 879 || pixel_index == 883 || pixel_index == 885 || pixel_index == 887 || pixel_index == 889 || pixel_index == 891 || pixel_index == 909 || pixel_index == 925 || pixel_index == 927 || pixel_index == 929 || pixel_index == 931 || pixel_index == 933 || pixel_index == 935 || pixel_index == 937 || pixel_index == 939 || pixel_index == 941 || pixel_index == 943 || pixel_index == 945 || pixel_index == 947 || pixel_index == 949 || pixel_index == 951 || pixel_index == 953 || pixel_index == 955 || pixel_index == 1061 || pixel_index == 1067 || pixel_index == 1073 || pixel_index == 1100 || pixel_index == 1117 || pixel_index == 1129 || pixel_index == 1135 || pixel_index == 1141 || pixel_index == 1147 || pixel_index == 1253 || pixel_index == 1309 || pixel_index == 1315 || pixel_index == 1317 || pixel_index == 1319 || pixel_index == 1321 || pixel_index == 1323 || pixel_index == 1325 || pixel_index == 1327 || pixel_index == 1329 || pixel_index == 1333 || pixel_index == 1335 || pixel_index == 1337 || pixel_index == 1339 || pixel_index == 1343 || pixel_index == 1389 || pixel_index == 1465 || pixel_index == 1508 || pixel_index == 1514 || pixel_index == 1520 || pixel_index == 1526 || pixel_index == 1565 || pixel_index == 1635 || pixel_index == 1657 || pixel_index == 1693 || pixel_index == 1715 || pixel_index == 1719 || pixel_index == 1721 || pixel_index == 1727 || pixel_index == 1843 || pixel_index == 1845 || pixel_index == 1885 || pixel_index == 1891 || pixel_index == 1901 || pixel_index == 1903 || pixel_index == 1909 || pixel_index == 1917 || pixel_index == 2019 || pixel_index == 2029 || pixel_index == 2031 || pixel_index == 2082 || pixel_index == 2084 || pixel_index == 2086 || pixel_index == 2104 || pixel_index == 2209 || pixel_index == 2223 || pixel_index == 2278 || pixel_index == 2286 || pixel_index == 2292 || pixel_index == 2302 || pixel_index == 2401 || pixel_index == 2403 || pixel_index == 2405 || pixel_index == 2413 || pixel_index == 2415 || pixel_index == 2417 || pixel_index == 2466 || pixel_index == 2468 || pixel_index == 2470 || pixel_index == 2478 || pixel_index == 2601 || pixel_index == 2613 || pixel_index == 2659 || pixel_index == 2785 || pixel_index == 2795 || pixel_index == 2859 || pixel_index == 2861 || pixel_index == 2867 || pixel_index == 2977 || pixel_index == 2991 || pixel_index == 2999 || pixel_index == 3050 || pixel_index == 3060 || pixel_index == 3062 || pixel_index == 3169 || pixel_index == 3177 || pixel_index == 3235 || pixel_index == 3352 || pixel_index == 3358 || pixel_index == 3367 || pixel_index == 3373 || pixel_index == 3379 || pixel_index == 3426 || pixel_index == 3436 || pixel_index == 3553 || pixel_index == 3619 || pixel_index == 3621 || pixel_index == 3734 || pixel_index == 3736 || pixel_index == 3745 || pixel_index == 3749 || pixel_index == 3761 || pixel_index == 3811 || pixel_index == 3928 || pixel_index == 3937 || pixel_index == 3945 || pixel_index == 3949 || pixel_index == 3951 || pixel_index == 3953 || pixel_index == 4008 || pixel_index == 4010 || pixel_index == 4145 || pixel_index == 4196 || pixel_index == 4200 || pixel_index == 4321 || pixel_index == 4327 || pixel_index == 4335 || pixel_index == 4341 || pixel_index == 4497 || pixel_index == 4513 || pixel_index == 4687 || pixel_index == 4689 || pixel_index == 4705 || pixel_index == 4717 || pixel_index == 4798 || pixel_index == 4880 || pixel_index == 4897 || pixel_index == 4901 || pixel_index == 4986 || pixel_index == 4988 || pixel_index == 4990 || pixel_index == 5267 || pixel_index == 5269 || pixel_index == 5479 || pixel_index == 5481 || pixel_index == 5483 || pixel_index == 5562 || pixel_index == 5673 || pixel_index == 5685 || pixel_index == 5688 || pixel_index == 5721 || pixel_index == 5830 || pixel_index == 5863 || pixel_index == 5865 || pixel_index == 5867 || pixel_index == 5869 || pixel_index == 5912 || pixel_index == 5914 || pixel_index == 5916 || pixel_index == 5930 || pixel_index == 5950 || pixel_index == 5992 || pixel_index == 6057 || pixel_index == 6108 || pixel_index == 6110 || pixel_index == 6126 || pixel_index == 6128 || pixel_index == 6130 || pixel_index == 6132) oled_data = 16'b0101101110010001;
    else if (pixel_index == 295 || pixel_index == 297 || pixel_index == 301 || pixel_index == 303 || pixel_index == 307 || pixel_index == 309 || pixel_index == 313 || pixel_index == 315 || pixel_index == 319 || pixel_index == 321 || pixel_index == 329 || pixel_index == 331 || pixel_index == 335 || pixel_index == 349 || pixel_index == 351 || pixel_index == 355 || pixel_index == 357 || pixel_index == 361 || pixel_index == 363 || pixel_index == 367 || pixel_index == 369 || pixel_index == 373 || pixel_index == 375 || pixel_index == 379 || pixel_index == 381 || pixel_index == 383 || pixel_index == 544 || pixel_index == 552 || pixel_index == 554 || pixel_index == 556 || pixel_index == 564 || pixel_index == 566 || pixel_index == 568 || pixel_index == 574 || pixel_index == 622 || pixel_index == 681 || pixel_index == 683 || pixel_index == 687 || pixel_index == 689 || pixel_index == 693 || pixel_index == 695 || pixel_index == 699 || pixel_index == 701 || pixel_index == 716 || pixel_index == 735 || pixel_index == 737 || pixel_index == 741 || pixel_index == 743 || pixel_index == 747 || pixel_index == 749 || pixel_index == 753 || pixel_index == 755 || pixel_index == 759 || pixel_index == 761 || pixel_index == 765 || pixel_index == 957 || pixel_index == 959 || pixel_index == 988 || pixel_index == 1063 || pixel_index == 1065 || pixel_index == 1069 || pixel_index == 1075 || pixel_index == 1083 || pixel_index == 1125 || pixel_index == 1127 || pixel_index == 1131 || pixel_index == 1133 || pixel_index == 1137 || pixel_index == 1139 || pixel_index == 1143 || pixel_index == 1145 || pixel_index == 1149 || pixel_index == 1151 || pixel_index == 1181 || pixel_index == 1198 || pixel_index == 1255 || pixel_index == 1265 || pixel_index == 1273 || pixel_index == 1275 || pixel_index == 1341 || pixel_index == 1373 || pixel_index == 1445 || pixel_index == 1447 || pixel_index == 1457 || pixel_index == 1467 || pixel_index == 1500 || pixel_index == 1506 || pixel_index == 1510 || pixel_index == 1512 || pixel_index == 1516 || pixel_index == 1518 || pixel_index == 1522 || pixel_index == 1524 || pixel_index == 1528 || pixel_index == 1532 || pixel_index == 1534 || pixel_index == 1637 || pixel_index == 1647 || pixel_index == 1659 || pixel_index == 1695 || pixel_index == 1697 || pixel_index == 1703 || pixel_index == 1705 || pixel_index == 1717 || pixel_index == 1723 || pixel_index == 1725 || pixel_index == 1758 || pixel_index == 1827 || pixel_index == 1839 || pixel_index == 1841 || pixel_index == 1847 || pixel_index == 1849 || pixel_index == 1889 || pixel_index == 1893 || pixel_index == 1895 || pixel_index == 1897 || pixel_index == 1899 || pixel_index == 1905 || pixel_index == 1907 || pixel_index == 1913 || pixel_index == 1915 || pixel_index == 1950 || pixel_index == 2027 || pixel_index == 2037 || pixel_index == 2039 || pixel_index == 2041 || pixel_index == 2076 || pixel_index == 2080 || pixel_index == 2088 || pixel_index == 2090 || pixel_index == 2092 || pixel_index == 2094 || pixel_index == 2096 || pixel_index == 2098 || pixel_index == 2100 || pixel_index == 2106 || pixel_index == 2108 || pixel_index == 2139 || pixel_index == 2141 || pixel_index == 2221 || pixel_index == 2225 || pixel_index == 2227 || pixel_index == 2229 || pixel_index == 2231 || pixel_index == 2233 || pixel_index == 2270 || pixel_index == 2272 || pixel_index == 2274 || pixel_index == 2276 || pixel_index == 2280 || pixel_index == 2282 || pixel_index == 2284 || pixel_index == 2288 || pixel_index == 2290 || pixel_index == 2296 || pixel_index == 2298 || pixel_index == 2300 || pixel_index == 2331 || pixel_index == 2389 || pixel_index == 2399 || pixel_index == 2407 || pixel_index == 2409 || pixel_index == 2411 || pixel_index == 2419 || pixel_index == 2421 || pixel_index == 2423 || pixel_index == 2425 || pixel_index == 2464 || pixel_index == 2472 || pixel_index == 2480 || pixel_index == 2482 || pixel_index == 2484 || pixel_index == 2487 || pixel_index == 2489 || pixel_index == 2491 || pixel_index == 2493 || pixel_index == 2590 || pixel_index == 2593 || pixel_index == 2603 || pixel_index == 2605 || pixel_index == 2611 || pixel_index == 2615 || pixel_index == 2657 || pixel_index == 2661 || pixel_index == 2663 || pixel_index == 2669 || pixel_index == 2671 || pixel_index == 2673 || pixel_index == 2675 || pixel_index == 2677 || pixel_index == 2679 || pixel_index == 2681 || pixel_index == 2683 || pixel_index == 2712 || pixel_index == 2780 || pixel_index == 2782 || pixel_index == 2791 || pixel_index == 2793 || pixel_index == 2803 || pixel_index == 2805 || pixel_index == 2807 || pixel_index == 2851 || pixel_index == 2853 || pixel_index == 2855 || pixel_index == 2857 || pixel_index == 2863 || pixel_index == 2865 || pixel_index == 2869 || pixel_index == 2871 || pixel_index == 2873 || pixel_index == 2970 || pixel_index == 2972 || pixel_index == 2974 || pixel_index == 2979 || pixel_index == 2981 || pixel_index == 2983 || pixel_index == 2985 || pixel_index == 2987 || pixel_index == 2989 || pixel_index == 2993 || pixel_index == 2995 || pixel_index == 2997 || pixel_index == 3042 || pixel_index == 3044 || pixel_index == 3048 || pixel_index == 3052 || pixel_index == 3054 || pixel_index == 3056 || pixel_index == 3058 || pixel_index == 3064 || pixel_index == 3162 || pixel_index == 3166 || pixel_index == 3173 || pixel_index == 3175 || pixel_index == 3179 || pixel_index == 3185 || pixel_index == 3187 || pixel_index == 3189 || pixel_index == 3239 || pixel_index == 3241 || pixel_index == 3243 || pixel_index == 3245 || pixel_index == 3247 || pixel_index == 3249 || pixel_index == 3251 || pixel_index == 3253 || pixel_index == 3255 || pixel_index == 3354 || pixel_index == 3356 || pixel_index == 3361 || pixel_index == 3363 || pixel_index == 3365 || pixel_index == 3371 || pixel_index == 3375 || pixel_index == 3377 || pixel_index == 3428 || pixel_index == 3430 || pixel_index == 3438 || pixel_index == 3440 || pixel_index == 3442 || pixel_index == 3444 || pixel_index == 3446 || pixel_index == 3543 || pixel_index == 3545 || pixel_index == 3549 || pixel_index == 3551 || pixel_index == 3555 || pixel_index == 3557 || pixel_index == 3559 || pixel_index == 3563 || pixel_index == 3565 || pixel_index == 3567 || pixel_index == 3569 || pixel_index == 3571 || pixel_index == 3573 || pixel_index == 3575 || pixel_index == 3623 || pixel_index == 3625 || pixel_index == 3627 || pixel_index == 3629 || pixel_index == 3631 || pixel_index == 3633 || pixel_index == 3635 || pixel_index == 3637 || pixel_index == 3738 || pixel_index == 3747 || pixel_index == 3759 || pixel_index == 3763 || pixel_index == 3765 || pixel_index == 3813 || pixel_index == 3815 || pixel_index == 3817 || pixel_index == 3819 || pixel_index == 3821 || pixel_index == 3823 || pixel_index == 3825 || pixel_index == 3827 || pixel_index == 3862 || pixel_index == 3906 || pixel_index == 3924 || pixel_index == 3926 || pixel_index == 3930 || pixel_index == 3932 || pixel_index == 3934 || pixel_index == 3939 || pixel_index == 3941 || pixel_index == 3943 || pixel_index == 3947 || pixel_index == 3960 || pixel_index == 4004 || pixel_index == 4006 || pixel_index == 4012 || pixel_index == 4014 || pixel_index == 4096 || pixel_index == 4098 || pixel_index == 4115 || pixel_index == 4117 || pixel_index == 4121 || pixel_index == 4123 || pixel_index == 4125 || pixel_index == 4127 || pixel_index == 4129 || pixel_index == 4131 || pixel_index == 4133 || pixel_index == 4135 || pixel_index == 4137 || pixel_index == 4139 || pixel_index == 4141 || pixel_index == 4143 || pixel_index == 4151 || pixel_index == 4198 || pixel_index == 4204 || pixel_index == 4206 || pixel_index == 4208 || pixel_index == 4305 || pixel_index == 4307 || pixel_index == 4309 || pixel_index == 4313 || pixel_index == 4315 || pixel_index == 4317 || pixel_index == 4323 || pixel_index == 4325 || pixel_index == 4329 || pixel_index == 4331 || pixel_index == 4333 || pixel_index == 4388 || pixel_index == 4390 || pixel_index == 4392 || pixel_index == 4394 || pixel_index == 4396 || pixel_index == 4398 || pixel_index == 4414 || pixel_index == 4495 || pixel_index == 4499 || pixel_index == 4507 || pixel_index == 4515 || pixel_index == 4517 || pixel_index == 4519 || pixel_index == 4521 || pixel_index == 4523 || pixel_index == 4525 || pixel_index == 4527 || pixel_index == 4583 || pixel_index == 4711 || pixel_index == 4778 || pixel_index == 4780 || pixel_index == 4794 || pixel_index == 4796 || pixel_index == 4878 || pixel_index == 4899 || pixel_index == 4903 || pixel_index == 4905 || pixel_index == 4907 || pixel_index == 5095 || pixel_index == 5097 || pixel_index == 5099 || pixel_index == 5103 || pixel_index == 5263 || pixel_index == 5265 || pixel_index == 5287 || pixel_index == 5293 || pixel_index == 5357 || pixel_index == 5366 || pixel_index == 5368 || pixel_index == 5370 || pixel_index == 5372 || pixel_index == 5374 || pixel_index == 5455 || pixel_index == 5457 || pixel_index == 5459 || pixel_index == 5475 || pixel_index == 5477 || pixel_index == 5545 || pixel_index == 5549 || pixel_index == 5556 || pixel_index == 5558 || pixel_index == 5560 || pixel_index == 5564 || pixel_index == 5566 || pixel_index == 5587 || pixel_index == 5590 || pixel_index == 5608 || pixel_index == 5612 || pixel_index == 5616 || pixel_index == 5619 || pixel_index == 5643 || pixel_index == 5669 || pixel_index == 5671 || pixel_index == 5675 || pixel_index == 5677 || pixel_index == 5679 || pixel_index == 5681 || pixel_index == 5690 || pixel_index == 5699 || pixel_index == 5701 || pixel_index == 5710 || pixel_index == 5714 || pixel_index == 5725 || pixel_index == 5727 || pixel_index == 5729 || pixel_index == 5731 || pixel_index == 5736 || pixel_index == 5746 || pixel_index == 5758 || pixel_index == 5779 || pixel_index == 5787 || pixel_index == 5798 || pixel_index == 5800 || pixel_index == 5804 || pixel_index == 5808 || pixel_index == 5828 || pixel_index == 5859 || pixel_index == 5861 || pixel_index == 5871 || pixel_index == 5873 || pixel_index == 5877 || pixel_index == 5879 || pixel_index == 5886 || pixel_index == 5888 || pixel_index == 5890 || pixel_index == 5918 || pixel_index == 5920 || pixel_index == 5922 || pixel_index == 5936 || pixel_index == 5948 || pixel_index == 5971 || pixel_index == 5979 || pixel_index == 5990 || pixel_index == 5996 || pixel_index == 6000 || pixel_index == 6027 || pixel_index == 6029 || pixel_index == 6051 || pixel_index == 6053 || pixel_index == 6055 || pixel_index == 6059 || pixel_index == 6061 || pixel_index == 6063 || pixel_index == 6071 || pixel_index == 6076 || pixel_index == 6078 || pixel_index == 6080 || pixel_index == 6082 || pixel_index == 6094 || pixel_index == 6098 || pixel_index == 6100 || pixel_index == 6102 || pixel_index == 6104 || pixel_index == 6106 || pixel_index == 6112 || pixel_index == 6114 || pixel_index == 6134 || pixel_index == 6136 || pixel_index == 6138 || pixel_index == 6140 || pixel_index == 6142) oled_data = 16'b0101001110010001;
    else if (pixel_index == 296 || pixel_index == 302 || pixel_index == 308 || pixel_index == 314 || pixel_index == 320 || pixel_index == 330 || pixel_index == 350 || pixel_index == 356 || pixel_index == 362 || pixel_index == 368 || pixel_index == 374 || pixel_index == 380 || pixel_index == 431 || pixel_index == 553 || pixel_index == 555 || pixel_index == 565 || pixel_index == 567 || pixel_index == 669 || pixel_index == 682 || pixel_index == 694 || pixel_index == 736 || pixel_index == 742 || pixel_index == 754 || pixel_index == 861 || pixel_index == 989 || pixel_index == 1102 || pixel_index == 1126 || pixel_index == 1132 || pixel_index == 1180 || pixel_index == 1245 || pixel_index == 1372 || pixel_index == 1437 || pixel_index == 1517 || pixel_index == 1563 || pixel_index == 1609 || pixel_index == 1621 || pixel_index == 1696 || pixel_index == 1742 || pixel_index == 1800 || pixel_index == 1840 || pixel_index == 1854 || pixel_index == 1984 || pixel_index == 1992 || pixel_index == 2001 || pixel_index == 2009 || pixel_index == 2011 || pixel_index == 2045 || pixel_index == 2091 || pixel_index == 2093 || pixel_index == 2176 || pixel_index == 2226 || pixel_index == 2235 || pixel_index == 2283 || pixel_index == 2324 || pixel_index == 2326 || pixel_index == 2376 || pixel_index == 2408 || pixel_index == 2494 || pixel_index == 2515 || pixel_index == 2560 || pixel_index == 2568 || pixel_index == 2585 || pixel_index == 2676 || pixel_index == 2700 || pixel_index == 2707 || pixel_index == 2808 || pixel_index == 2874 || pixel_index == 2900 || pixel_index == 2959 || pixel_index == 2961 || pixel_index == 2973 || pixel_index == 2980 || pixel_index == 3067 || pixel_index == 3071 || pixel_index == 3084 || pixel_index == 3092 || pixel_index == 3144 || pixel_index == 3242 || pixel_index == 3254 || pixel_index == 3335 || pixel_index == 3344 || pixel_index == 3429 || pixel_index == 3453 || pixel_index == 3467 || pixel_index == 3539 || pixel_index == 3558 || pixel_index == 3566 || pixel_index == 3642 || pixel_index == 3651 || pixel_index == 3729 || pixel_index == 3764 || pixel_index == 3843 || pixel_index == 3863 || pixel_index == 3916 || pixel_index == 3942 || pixel_index == 4001 || pixel_index == 4020 || pixel_index == 4022 || pixel_index == 4026 || pixel_index == 4036 || pixel_index == 4134 || pixel_index == 4136 || pixel_index == 4193 || pixel_index == 4213 || pixel_index == 4246 || pixel_index == 4413 || pixel_index == 4615 || pixel_index == 4680 || pixel_index == 4795 || pixel_index == 4812 || pixel_index == 4904 || pixel_index == 5003 || pixel_index == 5198 || pixel_index == 5369 || pixel_index == 5371 || pixel_index == 5373 || pixel_index == 5460 || pixel_index == 5476 || pixel_index == 5565 || pixel_index == 5586 || pixel_index == 5670 || pixel_index == 5676 || pixel_index == 5708 || pixel_index == 5726 || pixel_index == 5728 || pixel_index == 5732 || pixel_index == 5738 || pixel_index == 5876 || pixel_index == 5878 || pixel_index == 5919 || pixel_index == 5956 || pixel_index == 5968 || pixel_index == 6028 || pixel_index == 6054 || pixel_index == 6060 || pixel_index == 6093 || pixel_index == 6105 || pixel_index == 6115 || pixel_index == 6137 || pixel_index == 6141) oled_data = 16'b0101101101010010;
    else if (((pixel_index >= 435) && (pixel_index <= 438)) || ((pixel_index >= 516) && (pixel_index <= 518)) || ((pixel_index >= 531) && (pixel_index <= 535)) || ((pixel_index >= 611) && (pixel_index <= 615)) || ((pixel_index >= 626) && (pixel_index <= 631)) || ((pixel_index >= 706) && (pixel_index <= 712)) || ((pixel_index >= 721) && (pixel_index <= 723)) || ((pixel_index >= 727) && (pixel_index <= 728)) || ((pixel_index >= 801) && (pixel_index <= 803)) || ((pixel_index >= 806) && (pixel_index <= 808)) || ((pixel_index >= 817) && (pixel_index <= 818)) || ((pixel_index >= 823) && (pixel_index <= 824)) || ((pixel_index >= 897) && (pixel_index <= 899)) || ((pixel_index >= 903) && (pixel_index <= 904)) || ((pixel_index >= 913) && (pixel_index <= 914)) || ((pixel_index >= 919) && (pixel_index <= 921)) || ((pixel_index >= 993) && (pixel_index <= 994)) || ((pixel_index >= 999) && (pixel_index <= 1001)) || ((pixel_index >= 1009) && (pixel_index <= 1010)) || ((pixel_index >= 1015) && (pixel_index <= 1017)) || ((pixel_index >= 1088) && (pixel_index <= 1090)) || ((pixel_index >= 1096) && (pixel_index <= 1097)) || ((pixel_index >= 1105) && (pixel_index <= 1106)) || ((pixel_index >= 1112) && (pixel_index <= 1113)) || ((pixel_index >= 1184) && (pixel_index <= 1186)) || ((pixel_index >= 1192) && (pixel_index <= 1193)) || ((pixel_index >= 1201) && (pixel_index <= 1202)) || ((pixel_index >= 1208) && (pixel_index <= 1209)) || ((pixel_index >= 1281) && (pixel_index <= 1282)) || ((pixel_index >= 1288) && (pixel_index <= 1289)) || ((pixel_index >= 1297) && (pixel_index <= 1298)) || ((pixel_index >= 1304) && (pixel_index <= 1305)) || ((pixel_index >= 1377) && (pixel_index <= 1378)) || ((pixel_index >= 1384) && (pixel_index <= 1386)) || ((pixel_index >= 1393) && (pixel_index <= 1394)) || ((pixel_index >= 1400) && (pixel_index <= 1401)) || ((pixel_index >= 1473) && (pixel_index <= 1474)) || ((pixel_index >= 1480) && (pixel_index <= 1482)) || ((pixel_index >= 1489) && (pixel_index <= 1490)) || ((pixel_index >= 1496) && (pixel_index <= 1497)) || ((pixel_index >= 1569) && (pixel_index <= 1571)) || ((pixel_index >= 1577) && (pixel_index <= 1578)) || ((pixel_index >= 1585) && (pixel_index <= 1586)) || ((pixel_index >= 1592) && (pixel_index <= 1593)) || ((pixel_index >= 1665) && (pixel_index <= 1667)) || ((pixel_index >= 1673) && (pixel_index <= 1674)) || ((pixel_index >= 1681) && (pixel_index <= 1682)) || ((pixel_index >= 1688) && (pixel_index <= 1689)) || ((pixel_index >= 1762) && (pixel_index <= 1763)) || ((pixel_index >= 1769) && (pixel_index <= 1771)) || ((pixel_index >= 1777) && (pixel_index <= 1778)) || ((pixel_index >= 1783) && (pixel_index <= 1785)) || ((pixel_index >= 1858) && (pixel_index <= 1859)) || ((pixel_index >= 1865) && (pixel_index <= 1867)) || ((pixel_index >= 1874) && (pixel_index <= 1875)) || ((pixel_index >= 1879) && (pixel_index <= 1880)) || ((pixel_index >= 1954) && (pixel_index <= 1956)) || ((pixel_index >= 1961) && (pixel_index <= 1963)) || ((pixel_index >= 1970) && (pixel_index <= 1972)) || ((pixel_index >= 1974) && (pixel_index <= 1976)) || ((pixel_index >= 2051) && (pixel_index <= 2053)) || ((pixel_index >= 2056) && (pixel_index <= 2072)) || ((pixel_index >= 2147) && (pixel_index <= 2168)) || ((pixel_index >= 2243) && (pixel_index <= 2265)) || ((pixel_index >= 2336) && (pixel_index <= 2362)) || ((pixel_index >= 2430) && (pixel_index <= 2459)) || ((pixel_index >= 2525) && (pixel_index <= 2556)) || ((pixel_index >= 2621) && (pixel_index <= 2653)) || ((pixel_index >= 2716) && (pixel_index <= 2749)) || ((pixel_index >= 2812) && (pixel_index <= 2846)) || ((pixel_index >= 2907) && (pixel_index <= 2915)) || ((pixel_index >= 2921) && (pixel_index <= 2929)) || ((pixel_index >= 2935) && (pixel_index <= 2942)) || ((pixel_index >= 3003) && (pixel_index <= 3010)) || ((pixel_index >= 3018) && (pixel_index <= 3024)) || ((pixel_index >= 3032) && (pixel_index <= 3039)) || ((pixel_index >= 3098) && (pixel_index <= 3105)) || pixel_index == 3111 || ((pixel_index >= 3115) && (pixel_index <= 3119)) || ((pixel_index >= 3123) && (pixel_index <= 3125)) || ((pixel_index >= 3129) && (pixel_index <= 3135)) || ((pixel_index >= 3194) && (pixel_index <= 3200)) || ((pixel_index >= 3204) && (pixel_index <= 3208)) || ((pixel_index >= 3211) && (pixel_index <= 3215)) || ((pixel_index >= 3218) && (pixel_index <= 3222)) || ((pixel_index >= 3225) && (pixel_index <= 3231)) || ((pixel_index >= 3290) && (pixel_index <= 3327)) || ((pixel_index >= 3386) && (pixel_index <= 3423)) || ((pixel_index >= 3482) && (pixel_index <= 3485)) || ((pixel_index >= 3489) && (pixel_index <= 3510)) || ((pixel_index >= 3514) && (pixel_index <= 3519)) || ((pixel_index >= 3578) && (pixel_index <= 3581)) || ((pixel_index >= 3585) && (pixel_index <= 3592)) || ((pixel_index >= 3601) && (pixel_index <= 3606)) || ((pixel_index >= 3610) && (pixel_index <= 3615)) || ((pixel_index >= 3674) && (pixel_index <= 3688)) || ((pixel_index >= 3691) && (pixel_index <= 3694)) || ((pixel_index >= 3697) && (pixel_index <= 3711)) || ((pixel_index >= 3771) && (pixel_index <= 3785)) || ((pixel_index >= 3788) && (pixel_index <= 3789)) || ((pixel_index >= 3792) && (pixel_index <= 3806)) || ((pixel_index >= 3868) && (pixel_index <= 3881)) || ((pixel_index >= 3884) && (pixel_index <= 3885)) || ((pixel_index >= 3888) && (pixel_index <= 3901)) || ((pixel_index >= 3965) && (pixel_index <= 3978)) || ((pixel_index >= 3983) && (pixel_index <= 3996)) || ((pixel_index >= 4063) && (pixel_index <= 4091)) || ((pixel_index >= 4161) && (pixel_index <= 4184)) || ((pixel_index >= 4259) && (pixel_index <= 4279)) || ((pixel_index >= 4348) && (pixel_index <= 4349)) || pixel_index == 4381 || ((pixel_index >= 4443) && (pixel_index <= 4447)) || ((pixel_index >= 4474) && (pixel_index <= 4478)) || ((pixel_index >= 4538) && (pixel_index <= 4543)) || ((pixel_index >= 4570) && (pixel_index <= 4574)) || ((pixel_index >= 4634) && (pixel_index <= 4640)) || ((pixel_index >= 4666) && (pixel_index <= 4670)) || ((pixel_index >= 4730) && (pixel_index <= 4735)) || ((pixel_index >= 4763) && (pixel_index <= 4766)) || (pixel_index >= 4827) && (pixel_index <= 4830)) oled_data = 16'b1111111111111111;
    else if (pixel_index == 724 || pixel_index == 726 || pixel_index == 804 || pixel_index == 819 || pixel_index == 821 || pixel_index == 900 || pixel_index == 902 || pixel_index == 916 || pixel_index == 918 || pixel_index == 996 || pixel_index == 998 || pixel_index == 1011 || pixel_index == 1013 || pixel_index == 1091 || pixel_index == 1095 || pixel_index == 1110 || pixel_index == 1188 || pixel_index == 1190 || pixel_index == 1203 || pixel_index == 1205 || pixel_index == 1283 || pixel_index == 1285 || pixel_index == 1287 || pixel_index == 1299 || ((pixel_index >= 1301) && (pixel_index <= 1302)) || pixel_index == 1379 || pixel_index == 1381 || pixel_index == 1383 || pixel_index == 1396 || ((pixel_index >= 1398) && (pixel_index <= 1399)) || pixel_index == 1476 || pixel_index == 1478 || pixel_index == 1491 || pixel_index == 1574 || pixel_index == 1576 || pixel_index == 1588 || pixel_index == 1590 || pixel_index == 1668 || pixel_index == 1670 || pixel_index == 1672 || pixel_index == 1683 || pixel_index == 1685 || pixel_index == 1765 || pixel_index == 1767 || pixel_index == 1780 || pixel_index == 1860 || pixel_index == 1862 || pixel_index == 1876 || pixel_index == 1878 || pixel_index == 1959 || pixel_index == 2054 || pixel_index == 3486 || pixel_index == 3488 || pixel_index == 3511 || pixel_index == 3513 || pixel_index == 3583 || pixel_index == 3608) oled_data = 16'b1111110100110110;
    else if (pixel_index == 725 || pixel_index == 805 || pixel_index == 820 || pixel_index == 822 || pixel_index == 901 || pixel_index == 915 || pixel_index == 995 || pixel_index == 997 || pixel_index == 1012 || pixel_index == 1014 || pixel_index == 1092 || pixel_index == 1094 || pixel_index == 1107 || pixel_index == 1109 || pixel_index == 1187 || pixel_index == 1189 || pixel_index == 1204 || ((pixel_index >= 1206) && (pixel_index <= 1207)) || pixel_index == 1286 || pixel_index == 1380 || pixel_index == 1395 || pixel_index == 1397 || pixel_index == 1475 || pixel_index == 1477 || pixel_index == 1479 || pixel_index == 1492 || ((pixel_index >= 1494) && (pixel_index <= 1495)) || pixel_index == 1573 || pixel_index == 1587 || pixel_index == 1589 || pixel_index == 1669 || pixel_index == 1671 || ((pixel_index >= 1686) && (pixel_index <= 1687)) || pixel_index == 1764 || pixel_index == 1768 || pixel_index == 1779 || pixel_index == 1781 || pixel_index == 1861 || pixel_index == 1863 || pixel_index == 1877 || pixel_index == 1958 || pixel_index == 1960 || pixel_index == 2055 || pixel_index == 3487 || pixel_index == 3512 || pixel_index == 3582 || pixel_index == 3584 || pixel_index == 3607) oled_data = 16'b1111110100110101;
    else if (pixel_index == 917 || pixel_index == 1191 || pixel_index == 1284 || pixel_index == 1300 || pixel_index == 1303 || pixel_index == 1382 || pixel_index == 1575 || pixel_index == 1684 || pixel_index == 1766 || pixel_index == 3609) oled_data = 16'b1111110011110101;
    else if (pixel_index == 1093 || pixel_index == 1108 || pixel_index == 1111 || pixel_index == 1493 || pixel_index == 1572 || pixel_index == 1591 || pixel_index == 1782 || pixel_index == 1864 || pixel_index == 1957 || pixel_index == 1973) oled_data = 16'b1111110011110110;
    else if (pixel_index == 4627 || pixel_index == 4648 || pixel_index == 4656 || pixel_index == 4658 || pixel_index == 4673 || pixel_index == 4675 || pixel_index == 4722 || pixel_index == 4725 || pixel_index == 4739 || pixel_index == 4819 || pixel_index == 4917 || pixel_index == 4919 || pixel_index == 4931 || pixel_index == 4935 || pixel_index == 4937 || pixel_index == 4945 || pixel_index == 4953 || pixel_index == 4960 || pixel_index == 4962 || pixel_index == 4972 || pixel_index == 5025 || pixel_index == 5028 || pixel_index == 5051 || pixel_index == 5067 || pixel_index == 5070 || pixel_index == 5107 || pixel_index == 5205 || pixel_index == 5213 || pixel_index == 5215 || pixel_index == 5217 || pixel_index == 5219 || pixel_index == 5221 || pixel_index == 5223 || pixel_index == 5225 || pixel_index == 5227 || pixel_index == 5229 || pixel_index == 5231 || pixel_index == 5234 || pixel_index == 5236 || pixel_index == 5239 || pixel_index == 5245 || pixel_index == 5328 || pixel_index == 5333 || pixel_index == 5336 || pixel_index == 5340 || pixel_index == 5397 || pixel_index == 5412 || pixel_index == 5417 || pixel_index == 5427 || pixel_index == 5429 || pixel_index == 5439 || pixel_index == 5441 || pixel_index == 5443) oled_data = 16'b1110100100000101;
    else if (pixel_index == 4628 || pixel_index == 4630 || pixel_index == 4645 || pixel_index == 4651 || pixel_index == 4653 || pixel_index == 4661 || pixel_index == 4742 || pixel_index == 4745 || pixel_index == 4750 || pixel_index == 4752 || pixel_index == 4758 || pixel_index == 4771 || pixel_index == 4914 || pixel_index == 4940 || pixel_index == 4942 || pixel_index == 4947 || pixel_index == 4951 || pixel_index == 5011 || pixel_index == 5014 || pixel_index == 5031 || pixel_index == 5039 || pixel_index == 5041 || pixel_index == 5044 || pixel_index == 5046 || pixel_index == 5048 || pixel_index == 5053 || pixel_index == 5055 || pixel_index == 5203 || pixel_index == 5209 || pixel_index == 5211 || pixel_index == 5242 || pixel_index == 5248 || pixel_index == 5250 || pixel_index == 5303 || pixel_index == 5306 || pixel_index == 5320 || pixel_index == 5323 || pixel_index == 5338 || pixel_index == 5342 || pixel_index == 5400 || pixel_index == 5402 || pixel_index == 5405 || pixel_index == 5408 || pixel_index == 5410 || pixel_index == 5414 || pixel_index == 5423) oled_data = 16'b1110100100000100;
    else if (pixel_index == 4629 || pixel_index == 4644 || pixel_index == 4646 || pixel_index == 4650 || pixel_index == 4652 || pixel_index == 4654 || pixel_index == 4660 || pixel_index == 4662 || pixel_index == 4759 || pixel_index == 4939 || pixel_index == 4941 || pixel_index == 4943 || pixel_index == 4948 || pixel_index == 4950 || pixel_index == 5010 || pixel_index == 5012 || pixel_index == 5016 || pixel_index == 5045 || pixel_index == 5047 || pixel_index == 5054 || pixel_index == 5162 || pixel_index == 5164 || pixel_index == 5202 || pixel_index == 5210 || pixel_index == 5241 || pixel_index == 5247 || pixel_index == 5249 || pixel_index == 5302 || pixel_index == 5304 || pixel_index == 5307 || pixel_index == 5310 || pixel_index == 5318 || pixel_index == 5401 || pixel_index == 5404 || pixel_index == 5407 || pixel_index == 5409 || pixel_index == 5415 || pixel_index == 5419 || pixel_index == 5421 || pixel_index == 5425 || pixel_index == 5434 || pixel_index == 5437) oled_data = 16'b1110100011000101;
    else if (pixel_index == 4643 || pixel_index == 4647 || pixel_index == 4649 || pixel_index == 4655 || pixel_index == 4657 || pixel_index == 4659 || pixel_index == 4663 || pixel_index == 4674 || pixel_index == 4676 || ((pixel_index >= 4723) && (pixel_index <= 4724)) || pixel_index == 4726 || ((pixel_index >= 4740) && (pixel_index <= 4741)) || pixel_index == 4744 || pixel_index == 4746 || ((pixel_index >= 4748) && (pixel_index <= 4749)) || ((pixel_index >= 4753) && (pixel_index <= 4754)) || ((pixel_index >= 4756) && (pixel_index <= 4757)) || ((pixel_index >= 4769) && (pixel_index <= 4770)) || pixel_index == 4818 || pixel_index == 4916 || pixel_index == 4930 || pixel_index == 4932 || pixel_index == 4934 || pixel_index == 4936 || pixel_index == 4938 || pixel_index == 4944 || pixel_index == 4946 || pixel_index == 4959 || pixel_index == 4961 || ((pixel_index >= 4970) && (pixel_index <= 4971)) || pixel_index == 5013 || pixel_index == 5015 || pixel_index == 5024 || pixel_index == 5026 || ((pixel_index >= 5029) && (pixel_index <= 5030)) || pixel_index == 5033 || pixel_index == 5035 || pixel_index == 5037 || pixel_index == 5043 || ((pixel_index >= 5049) && (pixel_index <= 5050)) || pixel_index == 5052 || pixel_index == 5056 || pixel_index == 5058 || pixel_index == 5066 || ((pixel_index >= 5068) && (pixel_index <= 5069)) || pixel_index == 5106 || pixel_index == 5204 || pixel_index == 5206 || pixel_index == 5208 || pixel_index == 5212 || pixel_index == 5214 || pixel_index == 5216 || pixel_index == 5218 || pixel_index == 5220 || pixel_index == 5222 || pixel_index == 5224 || pixel_index == 5226 || pixel_index == 5228 || pixel_index == 5230 || ((pixel_index >= 5232) && (pixel_index <= 5233)) || pixel_index == 5235 || pixel_index == 5238 || pixel_index == 5244 || pixel_index == 5299 || pixel_index == 5301 || pixel_index == 5309 || ((pixel_index >= 5312) && (pixel_index <= 5313)) || ((pixel_index >= 5315) && (pixel_index <= 5316)) || pixel_index == 5321 || ((pixel_index >= 5324) && (pixel_index <= 5325)) || pixel_index == 5327 || pixel_index == 5329 || ((pixel_index >= 5331) && (pixel_index <= 5332)) || ((pixel_index >= 5334) && (pixel_index <= 5335)) || pixel_index == 5337 || pixel_index == 5339 || pixel_index == 5341 || pixel_index == 5343 || pixel_index == 5345 || pixel_index == 5396 || pixel_index == 5398 || pixel_index == 5403 || pixel_index == 5406 || pixel_index == 5411 || pixel_index == 5413 || pixel_index == 5416 || pixel_index == 5418 || pixel_index == 5422 || pixel_index == 5426 || pixel_index == 5430 || pixel_index == 5432 || pixel_index == 5435 || pixel_index == 5440 || pixel_index == 5442) oled_data = 16'b1110100011000100;
    else if (pixel_index == 4678 || ((pixel_index >= 4774) && (pixel_index <= 4775)) || pixel_index == 4869 || ((pixel_index >= 4871) && (pixel_index <= 4872)) || pixel_index == 4964 || ((pixel_index >= 4966) && (pixel_index <= 4967)) || ((pixel_index >= 5060) && (pixel_index <= 5062)) || pixel_index == 5064 || pixel_index == 5157 || ((pixel_index >= 5159) && (pixel_index <= 5160)) || ((pixel_index >= 5252) && (pixel_index <= 5255)) || pixel_index == 5349) oled_data = 16'b1001101011000111;
    else if (pixel_index == 4743 || pixel_index == 4751 || pixel_index == 5032 || pixel_index == 5040 || pixel_index == 5042 || pixel_index == 5057 || pixel_index == 5243 || pixel_index == 5322) oled_data = 16'b1110000011000101;
    else if (pixel_index == 4747 || pixel_index == 4755 || pixel_index == 4933 || pixel_index == 5036 || pixel_index == 5207 || pixel_index == 5300 || pixel_index == 5314 || pixel_index == 5326 || pixel_index == 5344 || pixel_index == 5431) oled_data = 16'b1110000100000101;
    else if (pixel_index == 4773 || pixel_index == 4870 || pixel_index == 4873 || pixel_index == 4965 || pixel_index == 4968 || pixel_index == 5063 || pixel_index == 5156 || pixel_index == 5158 || pixel_index == 5256 || pixel_index == 5348 || pixel_index == 5350) oled_data = 16'b1001101011001000;
    else if (pixel_index == 4915 || pixel_index == 4918 || pixel_index == 4952 || pixel_index == 5027 || pixel_index == 5038 || pixel_index == 5108 || pixel_index == 5237 || pixel_index == 5240 || pixel_index == 5246 || pixel_index == 5305 || pixel_index == 5319 || pixel_index == 5346 || pixel_index == 5399 || pixel_index == 5424 || pixel_index == 5428 || pixel_index == 5438) oled_data = 16'b1110000011000100;
    else if (pixel_index == 4949 || pixel_index == 5034 || pixel_index == 5163 || pixel_index == 5308 || pixel_index == 5311 || pixel_index == 5317 || pixel_index == 5330 || pixel_index == 5420 || pixel_index == 5433 || pixel_index == 5436) oled_data = 16'b1110000100000100;
    else oled_data = 0;



    end

endmodule
